
library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
-- read delay is 2 cycles

entity twiddleRom8192 is
	port(clk: in std_logic;
			romAddr: in unsigned(10-1 downto 0);
			romData: out std_logic_vector(30-1 downto 0)
			);
end entity;
architecture a of twiddleRom8192 is
	constant romDepthOrder: integer := 10;
	constant romDepth: integer := 2**romDepthOrder;
	constant romWidth: integer := 30;
	--ram
	type ram1t is array(0 to romDepth-1) of
		std_logic_vector(romWidth-1 downto 0);
	signal rom: ram1t;
	signal addr1: unsigned(romDepthOrder-1 downto 0) := (others=>'0');
	signal data0,data1: std_logic_vector(romWidth-1 downto 0) := (others=>'0');
begin
	addr1 <= romAddr when rising_edge(clk);
	data0 <= rom(to_integer(addr1));
	data1 <= data0 when rising_edge(clk);
	romData <= data1;
	rom <= (
"000000000011001111111111111111" , "000000000110010111111111111111" , "000000001001011111111111111111" , "000000001100101111111111111111" , "000000001111110111111111111111" , "000000010010111111111111111111" , "000000010110000111111111111111" , "000000011001001111111111111111" , "000000011100010111111111111111" , "000000011111011111111111111111"
, "000000100010100111111111111111" , "000000100101110111111111111111" , "000000101000111111111111111110" , "000000101100000111111111111110" , "000000101111001111111111111110" , "000000110010010111111111111110" , "000000110101011111111111111101" , "000000111000100111111111111101" , "000000111011110111111111111101" , "000000111110111111111111111100"
, "000001000010000111111111111100" , "000001000101001111111111111011" , "000001001000010111111111111011" , "000001001011011111111111111010" , "000001001110100111111111111010" , "000001010001101111111111111001" , "000001010100111111111111111001" , "000001011000000111111111111000" , "000001011011001111111111111000" , "000001011110010111111111110111"
, "000001100001011111111111110111" , "000001100100100111111111110110" , "000001100111101111111111110110" , "000001101010110111111111110101" , "000001101110000111111111110100" , "000001110001001111111111110100" , "000001110100010111111111110011" , "000001110111011111111111110010" , "000001111010100111111111110001" , "000001111101101111111111110001"
, "000010000000110111111111110000" , "000010000011111111111111101111" , "000010000111001111111111101110" , "000010001010010111111111101101" , "000010001101011111111111101100" , "000010010000100111111111101100" , "000010010011101111111111101011" , "000010010110110111111111101010" , "000010011001111111111111101001" , "000010011101000111111111101000"
, "000010100000001111111111100111" , "000010100011011111111111100110" , "000010100110100111111111100101" , "000010101001101111111111100100" , "000010101100110111111111100011" , "000010101111111111111111100010" , "000010110011000111111111100001" , "000010110110001111111111100000" , "000010111001010111111111011110" , "000010111100011111111111011101"
, "000010111111101111111111011100" , "000011000010110111111111011011" , "000011000101111111111111011010" , "000011001001000111111111011001" , "000011001100001111111111010111" , "000011001111010111111111010110" , "000011010010011111111111010101" , "000011010101100111111111010011" , "000011011000101111111111010010" , "000011011011110111111111010001"
, "000011011111000111111111001111" , "000011100010001111111111001110" , "000011100101010111111111001101" , "000011101000011111111111001011" , "000011101011100111111111001010" , "000011101110101111111111001000" , "000011110001110111111111000111" , "000011110100111111111111000101" , "000011111000000111111111000100" , "000011111011001111111111000010"
, "000011111110010111111111000001" , "000100000001100111111110111111" , "000100000100101111111110111110" , "000100000111110111111110111100" , "000100001010111111111110111010" , "000100001110000111111110111001" , "000100010001001111111110110111" , "000100010100010111111110110101" , "000100010111011111111110110100" , "000100011010100111111110110010"
, "000100011101101111111110110000" , "000100100000110111111110101110" , "000100100011111111111110101101" , "000100100111000111111110101011" , "000100101010001111111110101001" , "000100101101011111111110100111" , "000100110000100111111110100101" , "000100110011101111111110100011" , "000100110110110111111110100010" , "000100111001111111111110100000"
, "000100111101000111111110011110" , "000101000000001111111110011100" , "000101000011010111111110011010" , "000101000110011111111110011000" , "000101001001100111111110010110" , "000101001100101111111110010100" , "000101001111110111111110010010" , "000101010010111111111110010000" , "000101010110000111111110001110" , "000101011001001111111110001011"
, "000101011100010111111110001001" , "000101011111011111111110000111" , "000101100010100111111110000101" , "000101100101101111111110000011" , "000101101000111111111110000001" , "000101101100000111111101111110" , "000101101111001111111101111100" , "000101110010010111111101111010" , "000101110101011111111101111000" , "000101111000100111111101110101"
, "000101111011101111111101110011" , "000101111110110111111101110001" , "000110000001111111111101101110" , "000110000101000111111101101100" , "000110001000001111111101101010" , "000110001011010111111101100111" , "000110001110011111111101100101" , "000110010001100111111101100010" , "000110010100101111111101100000" , "000110010111110111111101011101"
, "000110011010111111111101011011" , "000110011110000111111101011000" , "000110100001001111111101010110" , "000110100100010111111101010011" , "000110100111011111111101010000" , "000110101010100111111101001110" , "000110101101101111111101001011" , "000110110000110111111101001001" , "000110110011111111111101000110" , "000110110111000111111101000011"
, "000110111010001111111101000001" , "000110111101010111111100111110" , "000111000000011111111100111011" , "000111000011100111111100111000" , "000111000110101111111100110110" , "000111001001110111111100110011" , "000111001100111111111100110000" , "000111010000000111111100101101" , "000111010011001111111100101010" , "000111010110010111111100100111"
, "000111011001011111111100100100" , "000111011100100111111100100010" , "000111011111100111111100011111" , "000111100010101111111100011100" , "000111100101110111111100011001" , "000111101000111111111100010110" , "000111101100000111111100010011" , "000111101111001111111100010000" , "000111110010010111111100001101" , "000111110101011111111100001010"
, "000111111000100111111100000110" , "000111111011101111111100000011" , "000111111110110111111100000000" , "001000000001111111111011111101" , "001000000101000111111011111010" , "001000001000001111111011110111" , "001000001011010111111011110100" , "001000001110011111111011110000" , "001000010001100111111011101101" , "001000010100100111111011101010"
, "001000010111101111111011100111" , "001000011010110111111011100011" , "001000011101111111111011100000" , "001000100001000111111011011101" , "001000100100001111111011011001" , "001000100111010111111011010110" , "001000101010011111111011010011" , "001000101101100111111011001111" , "001000110000101111111011001100" , "001000110011110111111011001000"
, "001000110110110111111011000101" , "001000111001111111111011000001" , "001000111101000111111010111110" , "001001000000001111111010111010" , "001001000011010111111010110111" , "001001000110011111111010110011" , "001001001001100111111010110000" , "001001001100101111111010101100" , "001001001111101111111010101000" , "001001010010110111111010100101"
, "001001010101111111111010100001" , "001001011001000111111010011101" , "001001011100001111111010011010" , "001001011111010111111010010110" , "001001100010011111111010010010" , "001001100101011111111010001110" , "001001101000100111111010001011" , "001001101011101111111010000111" , "001001101110110111111010000011" , "001001110001111111111001111111"
, "001001110101000111111001111011" , "001001111000001111111001111000" , "001001111011001111111001110100" , "001001111110010111111001110000" , "001010000001011111111001101100" , "001010000100100111111001101000" , "001010000111101111111001100100" , "001010001010101111111001100000" , "001010001101110111111001011100" , "001010010000111111111001011000"
, "001010010100000111111001010100" , "001010010111001111111001010000" , "001010011010001111111001001100" , "001010011101010111111001001000" , "001010100000011111111001000011" , "001010100011100111111000111111" , "001010100110101111111000111011" , "001010101001101111111000110111" , "001010101100110111111000110011" , "001010101111111111111000101111"
, "001010110011000111111000101010" , "001010110110001111111000100110" , "001010111001001111111000100010" , "001010111100010111111000011110" , "001010111111011111111000011001" , "001011000010100111111000010101" , "001011000101100111111000010001" , "001011001000101111111000001100" , "001011001011110111111000001000" , "001011001110111111111000000011"
, "001011010001111111110111111111" , "001011010101000111110111111011" , "001011011000001111110111110110" , "001011011011010111110111110010" , "001011011110010111110111101101" , "001011100001011111110111101001" , "001011100100100111110111100100" , "001011100111100111110111100000" , "001011101010101111110111011011" , "001011101101110111110111010110"
, "001011110000111111110111010010" , "001011110011111111110111001101" , "001011110111000111110111001001" , "001011111010001111110111000100" , "001011111101001111110110111111" , "001100000000010111110110111010" , "001100000011011111110110110110" , "001100000110011111110110110001" , "001100001001100111110110101100" , "001100001100101111110110100111"
, "001100001111101111110110100011" , "001100010010110111110110011110" , "001100010101111111110110011001" , "001100011000111111110110010100" , "001100011100000111110110001111" , "001100011111001111110110001010" , "001100100010001111110110000101" , "001100100101010111110110000001" , "001100101000011111110101111100" , "001100101011011111110101110111"
, "001100101110100111110101110010" , "001100110001101111110101101101" , "001100110100101111110101101000" , "001100110111110111110101100011" , "001100111010110111110101011101" , "001100111101111111110101011000" , "001101000001000111110101010011" , "001101000100000111110101001110" , "001101000111001111110101001001" , "001101001010001111110101000100"
, "001101001101010111110100111111" , "001101010000011111110100111010" , "001101010011011111110100110100" , "001101010110100111110100101111" , "001101011001100111110100101010" , "001101011100101111110100100101" , "001101011111110111110100011111" , "001101100010110111110100011010" , "001101100101111111110100010101" , "001101101000111111110100001111"
, "001101101100000111110100001010" , "001101101111000111110100000101" , "001101110010001111110011111111" , "001101110101001111110011111010" , "001101111000010111110011110100" , "001101111011010111110011101111" , "001101111110011111110011101001" , "001110000001100111110011100100" , "001110000100100111110011011110" , "001110000111101111110011011001"
, "001110001010101111110011010011" , "001110001101110111110011001110" , "001110010000110111110011001000" , "001110010011111111110011000010" , "001110010110111111110010111101" , "001110011010000111110010110111" , "001110011101000111110010110001" , "001110100000001111110010101100" , "001110100011001111110010100110" , "001110100110001111110010100000"
, "001110101001010111110010011011" , "001110101100010111110010010101" , "001110101111011111110010001111" , "001110110010011111110010001001" , "001110110101100111110010000011" , "001110111000100111110001111110" , "001110111011101111110001111000" , "001110111110101111110001110010" , "001111000001110111110001101100" , "001111000100110111110001100110"
, "001111000111110111110001100000" , "001111001010111111110001011010" , "001111001101111111110001010100" , "001111010001000111110001001110" , "001111010100000111110001001000" , "001111010111000111110001000010" , "001111011010001111110000111100" , "001111011101001111110000110110" , "001111100000010111110000110000" , "001111100011010111110000101010"
, "001111100110010111110000100100" , "001111101001011111110000011110" , "001111101100011111110000011000" , "001111101111011111110000010001" , "001111110010100111110000001011" , "001111110101100111110000000101" , "001111111000101111101111111111" , "001111111011101111101111111001" , "001111111110101111101111110010" , "010000000001110111101111101100"
, "010000000100110111101111100110" , "010000000111110111101111011111" , "010000001010111111101111011001" , "010000001101111111101111010011" , "010000010000111111101111001100" , "010000010011111111101111000110" , "010000010111000111101110111111" , "010000011010000111101110111001" , "010000011101000111101110110011" , "010000100000001111101110101100"
, "010000100011001111101110100110" , "010000100110001111101110011111" , "010000101001001111101110011001" , "010000101100010111101110010010" , "010000101111010111101110001011" , "010000110010010111101110000101" , "010000110101010111101101111110" , "010000111000011111101101111000" , "010000111011011111101101110001" , "010000111110011111101101101010"
, "010001000001011111101101100100" , "010001000100100111101101011101" , "010001000111100111101101010110" , "010001001010100111101101010000" , "010001001101100111101101001001" , "010001010000100111101101000010" , "010001010011101111101100111011" , "010001010110101111101100110100" , "010001011001101111101100101110" , "010001011100101111101100100111"
, "010001011111101111101100100000" , "010001100010110111101100011001" , "010001100101110111101100010010" , "010001101000110111101100001011" , "010001101011110111101100000100" , "010001101110110111101011111101" , "010001110001110111101011110110" , "010001110100111111101011101111" , "010001110111111111101011101000" , "010001111010111111101011100001"
, "010001111101111111101011011010" , "010010000000111111101011010011" , "010010000011111111101011001100" , "010010000110111111101011000101" , "010010001001111111101010111110" , "010010001100111111101010110111" , "010010010000000111101010110000" , "010010010011000111101010101000" , "010010010110000111101010100001" , "010010011001000111101010011010"
, "010010011100000111101010010011" , "010010011111000111101010001100" , "010010100010000111101010000100" , "010010100101000111101001111101" , "010010101000000111101001110110" , "010010101011000111101001101110" , "010010101110000111101001100111" , "010010110001000111101001100000" , "010010110100000111101001011000" , "010010110111000111101001010001"
, "010010111010000111101001001001" , "010010111101000111101001000010" , "010011000000000111101000111011" , "010011000011000111101000110011" , "010011000110000111101000101100" , "010011001001000111101000100100" , "010011001100000111101000011101" , "010011001111000111101000010101" , "010011010010000111101000001110" , "010011010101000111101000000110"
, "010011011000000111100111111110" , "010011011011000111100111110111" , "010011011110000111100111101111" , "010011100001000111100111100111" , "010011100100000111100111100000" , "010011100111000111100111011000" , "010011101010000111100111010000" , "010011101101000111100111001001" , "010011110000000111100111000001" , "010011110010111111100110111001"
, "010011110101111111100110110001" , "010011111000111111100110101010" , "010011111011111111100110100010" , "010011111110111111100110011010" , "010100000001111111100110010010" , "010100000100111111100110001010" , "010100000111111111100110000010" , "010100001010110111100101111010" , "010100001101110111100101110010" , "010100010000110111100101101010"
, "010100010011110111100101100010" , "010100010110110111100101011011" , "010100011001110111100101010011" , "010100011100101111100101001010" , "010100011111101111100101000010" , "010100100010101111100100111010" , "010100100101101111100100110010" , "010100101000101111100100101010" , "010100101011100111100100100010" , "010100101110100111100100011010"
, "010100110001100111100100010010" , "010100110100100111100100001010" , "010100110111100111100100000001" , "010100111010011111100011111001" , "010100111101011111100011110001" , "010101000000011111100011101001" , "010101000011011111100011100001" , "010101000110010111100011011000" , "010101001001010111100011010000" , "010101001100010111100011001000"
, "010101001111001111100010111111" , "010101010010001111100010110111" , "010101010101001111100010101111" , "010101011000001111100010100110" , "010101011011000111100010011110" , "010101011110000111100010010101" , "010101100001000111100010001101" , "010101100011111111100010000101" , "010101100110111111100001111100" , "010101101001111111100001110100"
, "010101101100110111100001101011" , "010101101111110111100001100011" , "010101110010101111100001011010" , "010101110101101111100001010001" , "010101111000101111100001001001" , "010101111011100111100001000000" , "010101111110100111100000111000" , "010110000001100111100000101111" , "010110000100011111100000100110" , "010110000111011111100000011110"
, "010110001010010111100000010101" , "010110001101010111100000001100" , "010110010000001111100000000011" , "010110010011001111011111111011" , "010110010110001111011111110010" , "010110011001000111011111101001" , "010110011100000111011111100000" , "010110011110111111011111011000" , "010110100001111111011111001111" , "010110100100110111011111000110"
, "010110100111110111011110111101" , "010110101010101111011110110100" , "010110101101101111011110101011" , "010110110000100111011110100010" , "010110110011100111011110011001" , "010110110110011111011110010000" , "010110111001011111011110000111" , "010110111100010111011101111110" , "010110111111010111011101110101" , "010111000010001111011101101100"
, "010111000101000111011101100011" , "010111001000000111011101011010" , "010111001010111111011101010001" , "010111001101111111011101001000" , "010111010000110111011100111111" , "010111010011110111011100110110" , "010111010110101111011100101101" , "010111011001100111011100100011" , "010111011100100111011100011010" , "010111011111011111011100010001"
, "010111100010011111011100001000" , "010111100101010111011011111110" , "010111101000001111011011110101" , "010111101011001111011011101100" , "010111101110000111011011100011" , "010111110000111111011011011001" , "010111110011111111011011010000" , "010111110110110111011011000111" , "010111111001101111011010111101" , "010111111100101111011010110100"
, "010111111111100111011010101010" , "011000000010011111011010100001" , "011000000101010111011010011000" , "011000001000010111011010001110" , "011000001011001111011010000101" , "011000001110000111011001111011" , "011000010001000111011001110010" , "011000010011111111011001101000" , "011000010110110111011001011110" , "011000011001101111011001010101"
, "011000011100101111011001001011" , "011000011111100111011001000010" , "011000100010011111011000111000" , "011000100101010111011000101110" , "011000101000001111011000100101" , "011000101011001111011000011011" , "011000101110000111011000010001" , "011000110000111111011000001000" , "011000110011110111010111111110" , "011000110110101111010111110100"
, "011000111001100111010111101010" , "011000111100100111010111100001" , "011000111111011111010111010111" , "011001000010010111010111001101" , "011001000101001111010111000011" , "011001001000000111010110111001" , "011001001010111111010110101111" , "011001001101110111010110100110" , "011001010000101111010110011100" , "011001010011101111010110010010"
, "011001010110100111010110001000" , "011001011001011111010101111110" , "011001011100010111010101110100" , "011001011111001111010101101010" , "011001100010000111010101100000" , "011001100100111111010101010110" , "011001100111110111010101001100" , "011001101010101111010101000010" , "011001101101100111010100111000" , "011001110000011111010100101101"
, "011001110011010111010100100011" , "011001110110001111010100011001" , "011001111001000111010100001111" , "011001111011111111010100000101" , "011001111110110111010011111011" , "011010000001101111010011110000" , "011010000100100111010011100110" , "011010000111011111010011011100" , "011010001010010111010011010010" , "011010001101001111010011000111"
, "011010010000000111010010111101" , "011010010010111111010010110011" , "011010010101101111010010101000" , "011010011000100111010010011110" , "011010011011011111010010010100" , "011010011110010111010010001001" , "011010100001001111010001111111" , "011010100100000111010001110101" , "011010100110111111010001101010" , "011010101001110111010001100000"
, "011010101100100111010001010101" , "011010101111011111010001001011" , "011010110010010111010001000000" , "011010110101001111010000110110" , "011010111000000111010000101011" , "011010111010111111010000100001" , "011010111101101111010000010110" , "011011000000100111010000001011" , "011011000011011111010000000001" , "011011000110010111001111110110"
, "011011001001000111001111101011" , "011011001011111111001111100001" , "011011001110110111001111010110" , "011011010001101111001111001011" , "011011010100011111001111000001" , "011011010111010111001110110110" , "011011011010001111001110101011" , "011011011101000111001110100000" , "011011011111110111001110010110" , "011011100010101111001110001011"
, "011011100101100111001110000000" , "011011101000010111001101110101" , "011011101011001111001101101010" , "011011101110000111001101011111" , "011011110000110111001101010101" , "011011110011101111001101001010" , "011011110110100111001100111111" , "011011111001010111001100110100" , "011011111100001111001100101001" , "011011111110111111001100011110"
, "011100000001110111001100010011" , "011100000100101111001100001000" , "011100000111011111001011111101" , "011100001010010111001011110010" , "011100001101000111001011100111" , "011100001111111111001011011100" , "011100010010101111001011010000" , "011100010101100111001011000101" , "011100011000010111001010111010" , "011100011011001111001010101111"
, "011100011110000111001010100100" , "011100100000110111001010011001" , "011100100011101111001010001101" , "011100100110011111001010000010" , "011100101001001111001001110111" , "011100101100000111001001101100" , "011100101110110111001001100000" , "011100110001101111001001010101" , "011100110100011111001001001010" , "011100110111010111001000111111"
, "011100111010000111001000110011" , "011100111100111111001000101000" , "011100111111101111001000011100" , "011101000010011111001000010001" , "011101000101010111001000000110" , "011101001000000111000111111010" , "011101001010111111000111101111" , "011101001101101111000111100011" , "011101010000011111000111011000" , "011101010011010111000111001100"
, "011101010110000111000111000001" , "011101011000110111000110110101" , "011101011011101111000110101010" , "011101011110011111000110011110" , "011101100001001111000110010011" , "011101100100000111000110000111" , "011101100110110111000101111011" , "011101101001100111000101110000" , "011101101100010111000101100100" , "011101101111001111000101011000"
, "011101110001111111000101001101" , "011101110100101111000101000001" , "011101110111011111000100110101" , "011101111010010111000100101010" , "011101111101000111000100011110" , "011101111111110111000100010010" , "011110000010100111000100000110" , "011110000101010111000011111010" , "011110001000001111000011101111" , "011110001010111111000011100011"
, "011110001101101111000011010111" , "011110010000011111000011001011" , "011110010011001111000010111111" , "011110010101111111000010110011" , "011110011000101111000010100111" , "011110011011100111000010011011" , "011110011110010111000010001111" , "011110100001000111000010000011" , "011110100011110111000001110111" , "011110100110100111000001101011"
, "011110101001010111000001011111" , "011110101100000111000001010011" , "011110101110110111000001000111" , "011110110001100111000000111011" , "011110110100010111000000101111" , "011110110111000111000000100011" , "011110111001110111000000010111" , "011110111100100111000000001011" , "011110111111010110111111111111" , "011111000010000110111111110010"
, "011111000100110110111111100110" , "011111000111100110111111011010" , "011111001010010110111111001110" , "011111001101000110111111000010" , "011111001111110110111110110101" , "011111010010100110111110101001" , "011111010101010110111110011101" , "011111011000000110111110010000" , "011111011010110110111110000100" , "011111011101100110111101111000"
, "011111100000001110111101101011" , "011111100010111110111101011111" , "011111100101101110111101010011" , "011111101000011110111101000110" , "011111101011001110111100111010" , "011111101101111110111100101101" , "011111110000101110111100100001" , "011111110011010110111100010100" , "011111110110000110111100001000" , "011111111000110110111011111011"
, "011111111011100110111011101111" , "011111111110001110111011100010" , "100000000000111110111011010110" , "100000000011101110111011001001" , "100000000110011110111010111101" , "100000001001000110111010110000" , "100000001011110110111010100011" , "100000001110100110111010010111" , "100000010001010110111010001010" , "100000010011111110111001111101"
, "100000010110101110111001110001" , "100000011001011110111001100100" , "100000011100000110111001010111" , "100000011110110110111001001010" , "100000100001100110111000111110" , "100000100100001110111000110001" , "100000100110111110111000100100" , "100000101001101110111000010111" , "100000101100010110111000001010" , "100000101111000110110111111110"
, "100000110001101110110111110001" , "100000110100011110110111100100" , "100000110111001110110111010111" , "100000111001110110110111001010" , "100000111100100110110110111101" , "100000111111001110110110110000" , "100001000001111110110110100011" , "100001000100100110110110010110" , "100001000111010110110110001001" , "100001001001111110110101111100"
, "100001001100101110110101101111" , "100001001111010110110101100010" , "100001010010000110110101010101" , "100001010100101110110101001000" , "100001010111011110110100111011" , "100001011010000110110100101110" , "100001011100110110110100100001" , "100001011111011110110100010100" , "100001100010000110110100000110" , "100001100100110110110011111001"
, "100001100111011110110011101100" , "100001101010001110110011011111" , "100001101100110110110011010010" , "100001101111011110110011000100" , "100001110010001110110010110111" , "100001110100110110110010101010" , "100001110111011110110010011101" , "100001111010001110110010001111" , "100001111100110110110010000010" , "100001111111011110110001110101"
, "100010000010001110110001100111" , "100010000100110110110001011010" , "100010000111011110110001001100" , "100010001010000110110000111111" , "100010001100110110110000110010" , "100010001111011110110000100100" , "100010010010000110110000010111" , "100010010100101110110000001001" , "100010010111010110101111111100" , "100010011010000110101111101110"
, "100010011100101110101111100001" , "100010011111010110101111010011" , "100010100001111110101111000110" , "100010100100100110101110111000" , "100010100111001110101110101010" , "100010101001111110101110011101" , "100010101100100110101110001111" , "100010101111001110101110000010" , "100010110001110110101101110100" , "100010110100011110101101100110"
, "100010110111000110101101011001" , "100010111001101110101101001011" , "100010111100010110101100111101" , "100010111110111110101100110000" , "100011000001100110101100100010" , "100011000100001110101100010100" , "100011000110110110101100000110" , "100011001001011110101011111000" , "100011001100000110101011101011" , "100011001110101110101011011101"
, "100011010001010110101011001111" , "100011010011111110101011000001" , "100011010110100110101010110011" , "100011011001001110101010100101" , "100011011011110110101010010111" , "100011011110011110101010001001" , "100011100001000110101001111100" , "100011100011101110101001101110" , "100011100110010110101001100000" , "100011101000111110101001010010"
, "100011101011100110101001000100" , "100011101110000110101000110110" , "100011110000101110101000101000" , "100011110011010110101000011010" , "100011110101111110101000001011" , "100011111000100110100111111101" , "100011111011001110100111101111" , "100011111101101110100111100001" , "100100000000010110100111010011" , "100100000010111110100111000101"
, "100100000101100110100110110111" , "100100001000000110100110101001" , "100100001010101110100110011010" , "100100001101010110100110001100" , "100100001111111110100101111110" , "100100010010011110100101110000" , "100100010101000110100101100001" , "100100010111101110100101010011" , "100100011010001110100101000101" , "100100011100110110100100110111"
, "100100011111011110100100101000" , "100100100001111110100100011010" , "100100100100100110100100001100" , "100100100111001110100011111101" , "100100101001101110100011101111" , "100100101100010110100011100000" , "100100101110110110100011010010" , "100100110001011110100011000100" , "100100110100000110100010110101" , "100100110110100110100010100111"
, "100100111001001110100010011000" , "100100111011101110100010001010" , "100100111110010110100001111011" , "100101000000110110100001101101" , "100101000011011110100001011110" , "100101000101111110100001010000" , "100101001000100110100001000001" , "100101001011000110100000110010" , "100101001101101110100000100100" , "100101010000001110100000010101"
, "100101010010101110100000000110" , "100101010101010110011111111000" , "100101010111110110011111101001" , "100101011010011110011111011010" , "100101011100111110011111001100" , "100101011111011110011110111101" , "100101100010000110011110101110" , "100101100100100110011110100000" , "100101100111000110011110010001" , "100101101001101110011110000010"
, "100101101100001110011101110011" , "100101101110101110011101100100" , "100101110001010110011101010110" , "100101110011110110011101000111" , "100101110110010110011100111000" , "100101111000111110011100101001" , "100101111011011110011100011010" , "100101111101111110011100001011" , "100110000000011110011011111100" , "100110000010111110011011101101"
, "100110000101100110011011011110" , "100110001000000110011011010000" , "100110001010100110011011000001" , "100110001101000110011010110010" , "100110001111100110011010100011" , "100110010010001110011010010011" , "100110010100101110011010000100" , "100110010111001110011001110101" , "100110011001101110011001100110" , "100110011100001110011001010111"
, "100110011110101110011001001000" , "100110100001001110011000111001" , "100110100011101110011000101010" , "100110100110001110011000011011" , "100110101000101110011000001100" , "100110101011001110010111111100" , "100110101101101110010111101101" , "100110110000001110010111011110" , "100110110010101110010111001111" , "100110110101001110010111000000"
, "100110110111101110010110110000" , "100110111010001110010110100001" , "100110111100101110010110010010" , "100110111111001110010110000010" , "100111000001101110010101110011" , "100111000100001110010101100100" , "100111000110101110010101010100" , "100111001001001110010101000101" , "100111001011101110010100110110" , "100111001110001110010100100110"
, "100111010000100110010100010111" , "100111010011000110010100000111" , "100111010101100110010011111000" , "100111011000000110010011101001" , "100111011010100110010011011001" , "100111011101000110010011001010" , "100111011111011110010010111010" , "100111100001111110010010101011" , "100111100100011110010010011011" , "100111100110111110010010001011"
, "100111101001010110010001111100" , "100111101011110110010001101100" , "100111101110010110010001011101" , "100111110000101110010001001101" , "100111110011001110010000111110" , "100111110101101110010000101110" , "100111111000000110010000011110" , "100111111010100110010000001111" , "100111111101000110001111111111" , "100111111111011110001111101111"
, "101000000001111110001111011111" , "101000000100011110001111010000" , "101000000110110110001111000000" , "101000001001010110001110110000" , "101000001011101110001110100000" , "101000001110001110001110010001" , "101000010000100110001110000001" , "101000010011000110001101110001" , "101000010101100110001101100001" , "101000010111111110001101010001"
, "101000011010011110001101000010" , "101000011100110110001100110010" , "101000011111001110001100100010" , "101000100001101110001100010010" , "101000100100000110001100000010" , "101000100110100110001011110010" , "101000101000111110001011100010" , "101000101011011110001011010010" , "101000101101110110001011000010" , "101000110000001110001010110010"
, "101000110010101110001010100010" , "101000110101000110001010010010" , "101000110111011110001010000010" , "101000111001111110001001110010" , "101000111100010110001001100010" , "101000111110101110001001010010" , "101001000001001110001001000010" , "101001000011100110001000110010" , "101001000101111110001000100001" , "101001001000011110001000010001"
, "101001001010110110001000000001" , "101001001101001110000111110001" , "101001001111100110000111100001" , "101001010010000110000111010001" , "101001010100011110000111000000" , "101001010110110110000110110000" , "101001011001001110000110100000" , "101001011011100110000110010000" , "101001011101111110000101111111" , "101001100000011110000101101111"
, "101001100010110110000101011111" , "101001100101001110000101001110" , "101001100111100110000100111110" , "101001101001111110000100101110" , "101001101100010110000100011101" , "101001101110101110000100001101" , "101001110001000110000011111101" , "101001110011011110000011101100" , "101001110101110110000011011100" , "101001111000001110000011001011"
, "101001111010100110000010111011" , "101001111100111110000010101010" , "101001111111010110000010011010" , "101010000001101110000010001001" , "101010000100000110000001111001" , "101010000110011110000001101000" , "101010001000110110000001011000" , "101010001011001110000001000111" , "101010001101100110000000110111" , "101010001111111110000000100110"
, "101010010010001110000000010110" , "101010010100100110000000000101" , "101010010110111101111111110100" , "101010011001010101111111100100" , "101010011011101101111111010011" , "101010011110000101111111000010" , "101010100000010101111110110010" , "101010100010101101111110100001" , "101010100101000101111110010000" , "101010100111011101111110000000"
, "101010101001110101111101101111" , "101010101100000101111101011110" , "101010101110011101111101001101" , "101010110000110101111100111100" , "101010110011000101111100101100" , "101010110101011101111100011011" , "101010110111110101111100001010" , "101010111010000101111011111001" , "101010111100011101111011101000" , "101010111110110101111011010111"
, "101011000001000101111011000111" , "101011000011011101111010110110" , "101011000101101101111010100101" , "101011001000000101111010010100" , "101011001010011101111010000011" , "101011001100101101111001110010" , "101011001111000101111001100001" , "101011010001010101111001010000" , "101011010011101101111000111111" , "101011010101111101111000101110"
, "101011011000010101111000011101" , "101011011010100101111000001100" , "101011011100111101110111111011" , "101011011111001101110111101010" , "101011100001100101110111011001" , "101011100011110101110111001000" , "101011100110000101110110110111" , "101011101000011101110110100101" , "101011101010101101110110010100" , "101011101100111101110110000011"
, "101011101111010101110101110010" , "101011110001100101110101100001" , "101011110011111101110101010000" , "101011110110001101110100111110" , "101011111000011101110100101101" , "101011111010101101110100011100" , "101011111101000101110100001011" , "101011111111010101110011111001" , "101100000001100101110011101000" , "101100000011110101110011010111"
, "101100000110001101110011000101" , "101100001000011101110010110100" , "101100001010101101110010100011" , "101100001100111101110010010001" , "101100001111001101110010000000" , "101100010001100101110001101111" , "101100010011110101110001011101" , "101100010110000101110001001100" , "101100011000010101110000111010" , "101100011010100101110000101001"
, "101100011100110101110000011000" , "101100011111000101110000000110" , "101100100001010101101111110101" , "101100100011100101101111100011" , "101100100101110101101111010010" , "101100101000000101101111000000" , "101100101010010101101110101111" , "101100101100100101101110011101" , "101100101110110101101110001100" , "101100110001000101101101111010"
, "101100110011010101101101101000" , "101100110101100101101101010111" , "101100110111110101101101000101" , "101100111010000101101100110100" , "101100111100010101101100100010" , "101100111110100101101100010000" , "101101000000110101101011111111" , "101101000011000101101011101101" , "101101000101001101101011011011" , "101101000111011101101011001001"
, "101101001001101101101010111000" , "101101001011111101101010100110" , "101101001110001101101010010100" , "101101010000010101101010000010"
);
end a;

