
library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
-- read delay is 2 cycles

entity twiddleRom32768 is
	port(clk: in std_logic;
			romAddr: in unsigned(12-1 downto 0);
			romData: out std_logic_vector(30-1 downto 0)
			);
end entity;
architecture a of twiddleRom32768 is
	constant romDepthOrder: integer := 12;
	constant romDepth: integer := 2**romDepthOrder;
	constant romWidth: integer := 30;
	--ram
	type ram1t is array(0 to romDepth-1) of
		std_logic_vector(romWidth-1 downto 0);
	signal rom: ram1t;
	signal addr1: unsigned(romDepthOrder-1 downto 0) := (others=>'0');
	signal data0,data1: std_logic_vector(romWidth-1 downto 0) := (others=>'0');
begin
	addr1 <= romAddr when rising_edge(clk);
	data0 <= rom(to_integer(addr1));
	data1 <= data0 when rising_edge(clk);
	romData <= data1;
	rom <= (
"000000000000110111111111111111" , "000000000001101111111111111111" , "000000000010011111111111111111" , "000000000011001111111111111111" , "000000000011111111111111111111" , "000000000100110111111111111111" , "000000000101100111111111111111" , "000000000110010111111111111111" , "000000000111001111111111111111" , "000000000111111111111111111111"
, "000000001000101111111111111111" , "000000001001011111111111111111" , "000000001010010111111111111111" , "000000001011000111111111111111" , "000000001011110111111111111111" , "000000001100101111111111111111" , "000000001101011111111111111111" , "000000001110001111111111111111" , "000000001110111111111111111111" , "000000001111110111111111111111"
, "000000010000100111111111111111" , "000000010001010111111111111111" , "000000010010001111111111111111" , "000000010010111111111111111111" , "000000010011101111111111111111" , "000000010100011111111111111111" , "000000010101010111111111111111" , "000000010110000111111111111111" , "000000010110110111111111111111" , "000000010111100111111111111111"
, "000000011000011111111111111111" , "000000011001001111111111111111" , "000000011001111111111111111111" , "000000011010110111111111111111" , "000000011011100111111111111111" , "000000011100010111111111111111" , "000000011101000111111111111111" , "000000011101111111111111111111" , "000000011110101111111111111111" , "000000011111011111111111111111"
, "000000100000010111111111111111" , "000000100001000111111111111111" , "000000100001110111111111111111" , "000000100010100111111111111111" , "000000100011011111111111111111" , "000000100100001111111111111111" , "000000100100111111111111111111" , "000000100101110111111111111111" , "000000100110100111111111111111" , "000000100111010111111111111110"
, "000000101000000111111111111110" , "000000101000111111111111111110" , "000000101001101111111111111110" , "000000101010011111111111111110" , "000000101011010111111111111110" , "000000101100000111111111111110" , "000000101100110111111111111110" , "000000101101100111111111111110" , "000000101110011111111111111110" , "000000101111001111111111111110"
, "000000101111111111111111111110" , "000000110000110111111111111110" , "000000110001100111111111111110" , "000000110010010111111111111110" , "000000110011000111111111111101" , "000000110011111111111111111101" , "000000110100101111111111111101" , "000000110101011111111111111101" , "000000110110010111111111111101" , "000000110111000111111111111101"
, "000000110111110111111111111101" , "000000111000100111111111111101" , "000000111001011111111111111101" , "000000111010001111111111111101" , "000000111010111111111111111101" , "000000111011110111111111111101" , "000000111100100111111111111100" , "000000111101010111111111111100" , "000000111110000111111111111100" , "000000111110111111111111111100"
, "000000111111101111111111111100" , "000001000000011111111111111100" , "000001000001001111111111111100" , "000001000010000111111111111100" , "000001000010110111111111111100" , "000001000011100111111111111100" , "000001000100011111111111111011" , "000001000101001111111111111011" , "000001000101111111111111111011" , "000001000110101111111111111011"
, "000001000111100111111111111011" , "000001001000010111111111111011" , "000001001001000111111111111011" , "000001001001111111111111111011" , "000001001010101111111111111011" , "000001001011011111111111111010" , "000001001100001111111111111010" , "000001001101000111111111111010" , "000001001101110111111111111010" , "000001001110100111111111111010"
, "000001001111011111111111111010" , "000001010000001111111111111010" , "000001010000111111111111111010" , "000001010001101111111111111001" , "000001010010100111111111111001" , "000001010011010111111111111001" , "000001010100000111111111111001" , "000001010100111111111111111001" , "000001010101101111111111111001" , "000001010110011111111111111001"
, "000001010111001111111111111001" , "000001011000000111111111111000" , "000001011000110111111111111000" , "000001011001100111111111111000" , "000001011010011111111111111000" , "000001011011001111111111111000" , "000001011011111111111111111000" , "000001011100101111111111111000" , "000001011101100111111111110111" , "000001011110010111111111110111"
, "000001011111000111111111110111" , "000001011111110111111111110111" , "000001100000101111111111110111" , "000001100001011111111111110111" , "000001100010001111111111110111" , "000001100011000111111111110110" , "000001100011110111111111110110" , "000001100100100111111111110110" , "000001100101010111111111110110" , "000001100110001111111111110110"
, "000001100110111111111111110110" , "000001100111101111111111110110" , "000001101000100111111111110101" , "000001101001010111111111110101" , "000001101010000111111111110101" , "000001101010110111111111110101" , "000001101011101111111111110101" , "000001101100011111111111110101" , "000001101101001111111111110100" , "000001101110000111111111110100"
, "000001101110110111111111110100" , "000001101111100111111111110100" , "000001110000010111111111110100" , "000001110001001111111111110100" , "000001110001111111111111110011" , "000001110010101111111111110011" , "000001110011100111111111110011" , "000001110100010111111111110011" , "000001110101000111111111110011" , "000001110101110111111111110010"
, "000001110110101111111111110010" , "000001110111011111111111110010" , "000001111000001111111111110010" , "000001111000111111111111110010" , "000001111001110111111111110010" , "000001111010100111111111110001" , "000001111011010111111111110001" , "000001111100001111111111110001" , "000001111100111111111111110001" , "000001111101101111111111110001"
, "000001111110011111111111110000" , "000001111111010111111111110000" , "000010000000000111111111110000" , "000010000000110111111111110000" , "000010000001101111111111110000" , "000010000010011111111111101111" , "000010000011001111111111101111" , "000010000011111111111111101111" , "000010000100110111111111101111" , "000010000101100111111111101111"
, "000010000110010111111111101110" , "000010000111001111111111101110" , "000010000111111111111111101110" , "000010001000101111111111101110" , "000010001001011111111111101110" , "000010001010010111111111101101" , "000010001011000111111111101101" , "000010001011110111111111101101" , "000010001100100111111111101101" , "000010001101011111111111101100"
, "000010001110001111111111101100" , "000010001110111111111111101100" , "000010001111110111111111101100" , "000010010000100111111111101100" , "000010010001010111111111101011" , "000010010010000111111111101011" , "000010010010111111111111101011" , "000010010011101111111111101011" , "000010010100011111111111101010" , "000010010101010111111111101010"
, "000010010110000111111111101010" , "000010010110110111111111101010" , "000010010111100111111111101010" , "000010011000011111111111101001" , "000010011001001111111111101001" , "000010011001111111111111101001" , "000010011010101111111111101001" , "000010011011100111111111101000" , "000010011100010111111111101000" , "000010011101000111111111101000"
, "000010011101111111111111101000" , "000010011110101111111111100111" , "000010011111011111111111100111" , "000010100000001111111111100111" , "000010100001000111111111100111" , "000010100001110111111111100110" , "000010100010100111111111100110" , "000010100011011111111111100110" , "000010100100001111111111100110" , "000010100100111111111111100101"
, "000010100101101111111111100101" , "000010100110100111111111100101" , "000010100111010111111111100101" , "000010101000000111111111100100" , "000010101000111111111111100100" , "000010101001101111111111100100" , "000010101010011111111111100100" , "000010101011001111111111100011" , "000010101100000111111111100011" , "000010101100110111111111100011"
, "000010101101100111111111100011" , "000010101110010111111111100010" , "000010101111001111111111100010" , "000010101111111111111111100010" , "000010110000101111111111100010" , "000010110001100111111111100001" , "000010110010010111111111100001" , "000010110011000111111111100001" , "000010110011110111111111100000" , "000010110100101111111111100000"
, "000010110101011111111111100000" , "000010110110001111111111100000" , "000010110110111111111111011111" , "000010110111110111111111011111" , "000010111000100111111111011111" , "000010111001010111111111011110" , "000010111010001111111111011110" , "000010111010111111111111011110" , "000010111011101111111111011110" , "000010111100011111111111011101"
, "000010111101010111111111011101" , "000010111110000111111111011101" , "000010111110110111111111011100" , "000010111111101111111111011100" , "000011000000011111111111011100" , "000011000001001111111111011100" , "000011000001111111111111011011" , "000011000010110111111111011011" , "000011000011100111111111011011" , "000011000100010111111111011010"
, "000011000101000111111111011010" , "000011000101111111111111011010" , "000011000110101111111111011001" , "000011000111011111111111011001" , "000011001000010111111111011001" , "000011001001000111111111011001" , "000011001001110111111111011000" , "000011001010100111111111011000" , "000011001011011111111111011000" , "000011001100001111111111010111"
, "000011001100111111111111010111" , "000011001101110111111111010111" , "000011001110100111111111010110" , "000011001111010111111111010110" , "000011010000000111111111010110" , "000011010000111111111111010101" , "000011010001101111111111010101" , "000011010010011111111111010101" , "000011010011001111111111010100" , "000011010100000111111111010100"
, "000011010100110111111111010100" , "000011010101100111111111010011" , "000011010110011111111111010011" , "000011010111001111111111010011" , "000011010111111111111111010010" , "000011011000101111111111010010" , "000011011001100111111111010010" , "000011011010010111111111010001" , "000011011011000111111111010001" , "000011011011110111111111010001"
, "000011011100101111111111010000" , "000011011101011111111111010000" , "000011011110001111111111010000" , "000011011111000111111111001111" , "000011011111110111111111001111" , "000011100000100111111111001111" , "000011100001010111111111001110" , "000011100010001111111111001110" , "000011100010111111111111001110" , "000011100011101111111111001101"
, "000011100100011111111111001101" , "000011100101010111111111001101" , "000011100110000111111111001100" , "000011100110110111111111001100" , "000011100111101111111111001100" , "000011101000011111111111001011" , "000011101001001111111111001011" , "000011101001111111111111001011" , "000011101010110111111111001010" , "000011101011100111111111001010"
, "000011101100010111111111001001" , "000011101101000111111111001001" , "000011101101111111111111001001" , "000011101110101111111111001000" , "000011101111011111111111001000" , "000011110000010111111111001000" , "000011110001000111111111000111" , "000011110001110111111111000111" , "000011110010100111111111000110" , "000011110011011111111111000110"
, "000011110100001111111111000110" , "000011110100111111111111000101" , "000011110101101111111111000101" , "000011110110100111111111000101" , "000011110111010111111111000100" , "000011111000000111111111000100" , "000011111000111111111111000011" , "000011111001101111111111000011" , "000011111010011111111111000011" , "000011111011001111111111000010"
, "000011111100000111111111000010" , "000011111100110111111111000010" , "000011111101100111111111000001" , "000011111110010111111111000001" , "000011111111001111111111000000" , "000011111111111111111111000000" , "000100000000101111111111000000" , "000100000001100111111110111111" , "000100000010010111111110111111" , "000100000011000111111110111110"
, "000100000011110111111110111110" , "000100000100101111111110111110" , "000100000101011111111110111101" , "000100000110001111111110111101" , "000100000110111111111110111100" , "000100000111110111111110111100" , "000100001000100111111110111100" , "000100001001010111111110111011" , "000100001010001111111110111011" , "000100001010111111111110111010"
, "000100001011101111111110111010" , "000100001100011111111110111010" , "000100001101010111111110111001" , "000100001110000111111110111001" , "000100001110110111111110111000" , "000100001111100111111110111000" , "000100010000011111111110110111" , "000100010001001111111110110111" , "000100010001111111111110110111" , "000100010010101111111110110110"
, "000100010011100111111110110110" , "000100010100010111111110110101" , "000100010101000111111110110101" , "000100010101111111111110110101" , "000100010110101111111110110100" , "000100010111011111111110110100" , "000100011000001111111110110011" , "000100011001000111111110110011" , "000100011001110111111110110010" , "000100011010100111111110110010"
, "000100011011010111111110110010" , "000100011100001111111110110001" , "000100011100111111111110110001" , "000100011101101111111110110000" , "000100011110011111111110110000" , "000100011111010111111110101111" , "000100100000000111111110101111" , "000100100000110111111110101110" , "000100100001101111111110101110" , "000100100010011111111110101110"
, "000100100011001111111110101101" , "000100100011111111111110101101" , "000100100100110111111110101100" , "000100100101100111111110101100" , "000100100110010111111110101011" , "000100100111000111111110101011" , "000100100111111111111110101010" , "000100101000101111111110101010" , "000100101001011111111110101010" , "000100101010001111111110101001"
, "000100101011000111111110101001" , "000100101011110111111110101000" , "000100101100100111111110101000" , "000100101101011111111110100111" , "000100101110001111111110100111" , "000100101110111111111110100110" , "000100101111101111111110100110" , "000100110000100111111110100101" , "000100110001010111111110100101" , "000100110010000111111110100100"
, "000100110010110111111110100100" , "000100110011101111111110100011" , "000100110100011111111110100011" , "000100110101001111111110100011" , "000100110101111111111110100010" , "000100110110110111111110100010" , "000100110111100111111110100001" , "000100111000010111111110100001" , "000100111001001111111110100000" , "000100111001111111111110100000"
, "000100111010101111111110011111" , "000100111011011111111110011111" , "000100111100010111111110011110" , "000100111101000111111110011110" , "000100111101110111111110011101" , "000100111110100111111110011101" , "000100111111011111111110011100" , "000101000000001111111110011100" , "000101000000111111111110011011" , "000101000001101111111110011011"
, "000101000010100111111110011010" , "000101000011010111111110011010" , "000101000100000111111110011001" , "000101000100111111111110011001" , "000101000101101111111110011000" , "000101000110011111111110011000" , "000101000111001111111110010111" , "000101001000000111111110010111" , "000101001000110111111110010110" , "000101001001100111111110010110"
, "000101001010010111111110010101" , "000101001011001111111110010101" , "000101001011111111111110010100" , "000101001100101111111110010100" , "000101001101011111111110010011" , "000101001110010111111110010011" , "000101001111000111111110010010" , "000101001111110111111110010010" , "000101010000100111111110010001" , "000101010001011111111110010001"
, "000101010010001111111110010000" , "000101010010111111111110010000" , "000101010011101111111110001111" , "000101010100100111111110001111" , "000101010101010111111110001110" , "000101010110000111111110001110" , "000101010110111111111110001101" , "000101010111101111111110001101" , "000101011000011111111110001100" , "000101011001001111111110001011"
, "000101011010000111111110001011" , "000101011010110111111110001010" , "000101011011100111111110001010" , "000101011100010111111110001001" , "000101011101001111111110001001" , "000101011101111111111110001000" , "000101011110101111111110001000" , "000101011111011111111110000111" , "000101100000010111111110000111" , "000101100001000111111110000110"
, "000101100001110111111110000110" , "000101100010100111111110000101" , "000101100011011111111110000100" , "000101100100001111111110000100" , "000101100100111111111110000011" , "000101100101101111111110000011" , "000101100110100111111110000010" , "000101100111010111111110000010" , "000101101000000111111110000001" , "000101101000111111111110000001"
, "000101101001101111111110000000" , "000101101010011111111110000000" , "000101101011001111111101111111" , "000101101100000111111101111110" , "000101101100110111111101111110" , "000101101101100111111101111101" , "000101101110010111111101111101" , "000101101111001111111101111100" , "000101101111111111111101111100" , "000101110000101111111101111011"
, "000101110001011111111101111010" , "000101110010010111111101111010" , "000101110011000111111101111001" , "000101110011110111111101111001" , "000101110100100111111101111000" , "000101110101011111111101111000" , "000101110110001111111101110111" , "000101110110111111111101110110" , "000101110111101111111101110110" , "000101111000100111111101110101"
, "000101111001010111111101110101" , "000101111010000111111101110100" , "000101111010110111111101110100" , "000101111011101111111101110011" , "000101111100011111111101110010" , "000101111101001111111101110010" , "000101111101111111111101110001" , "000101111110110111111101110001" , "000101111111100111111101110000" , "000110000000010111111101101111"
, "000110000001000111111101101111" , "000110000001111111111101101110" , "000110000010101111111101101110" , "000110000011011111111101101101" , "000110000100010111111101101101" , "000110000101000111111101101100" , "000110000101110111111101101011" , "000110000110100111111101101011" , "000110000111011111111101101010" , "000110001000001111111101101010"
, "000110001000111111111101101001" , "000110001001101111111101101000" , "000110001010100111111101101000" , "000110001011010111111101100111" , "000110001100000111111101100110" , "000110001100110111111101100110" , "000110001101101111111101100101" , "000110001110011111111101100101" , "000110001111001111111101100100" , "000110001111111111111101100011"
, "000110010000110111111101100011" , "000110010001100111111101100010" , "000110010010010111111101100010" , "000110010011000111111101100001" , "000110010011111111111101100000" , "000110010100101111111101100000" , "000110010101011111111101011111" , "000110010110001111111101011110" , "000110010111000111111101011110" , "000110010111110111111101011101"
, "000110011000100111111101011101" , "000110011001010111111101011100" , "000110011010001111111101011011" , "000110011010111111111101011011" , "000110011011101111111101011010" , "000110011100011111111101011001" , "000110011101010111111101011001" , "000110011110000111111101011000" , "000110011110110111111101011000" , "000110011111100111111101010111"
, "000110100000011111111101010110" , "000110100001001111111101010110" , "000110100001111111111101010101" , "000110100010101111111101010100" , "000110100011100111111101010100" , "000110100100010111111101010011" , "000110100101000111111101010010" , "000110100101110111111101010010" , "000110100110101111111101010001" , "000110100111011111111101010000"
, "000110101000001111111101010000" , "000110101000111111111101001111" , "000110101001110111111101001111" , "000110101010100111111101001110" , "000110101011010111111101001101" , "000110101100000111111101001101" , "000110101100111111111101001100" , "000110101101101111111101001011" , "000110101110011111111101001011" , "000110101111001111111101001010"
, "000110110000000111111101001001" , "000110110000110111111101001001" , "000110110001100111111101001000" , "000110110010010111111101000111" , "000110110011001111111101000111" , "000110110011111111111101000110" , "000110110100101111111101000101" , "000110110101011111111101000101" , "000110110110010111111101000100" , "000110110111000111111101000011"
, "000110110111110111111101000011" , "000110111000100111111101000010" , "000110111001011111111101000001" , "000110111010001111111101000001" , "000110111010111111111101000000" , "000110111011101111111100111111" , "000110111100100111111100111111" , "000110111101010111111100111110" , "000110111110000111111100111101" , "000110111110110111111100111100"
, "000110111111101111111100111100" , "000111000000011111111100111011" , "000111000001001111111100111010" , "000111000001111111111100111010" , "000111000010110111111100111001" , "000111000011100111111100111000" , "000111000100010111111100111000" , "000111000101000111111100110111" , "000111000101110111111100110110" , "000111000110101111111100110110"
, "000111000111011111111100110101" , "000111001000001111111100110100" , "000111001000111111111100110011" , "000111001001110111111100110011" , "000111001010100111111100110010" , "000111001011010111111100110001" , "000111001100000111111100110001" , "000111001100111111111100110000" , "000111001101101111111100101111" , "000111001110011111111100101111"
, "000111001111001111111100101110" , "000111010000000111111100101101" , "000111010000110111111100101100" , "000111010001100111111100101100" , "000111010010010111111100101011" , "000111010011001111111100101010" , "000111010011111111111100101010" , "000111010100101111111100101001" , "000111010101011111111100101000" , "000111010110010111111100100111"
, "000111010111000111111100100111" , "000111010111110111111100100110" , "000111011000100111111100100101" , "000111011001011111111100100100" , "000111011010001111111100100100" , "000111011010111111111100100011" , "000111011011101111111100100010" , "000111011100100111111100100010" , "000111011101010111111100100001" , "000111011110000111111100100000"
, "000111011110110111111100011111" , "000111011111100111111100011111" , "000111100000011111111100011110" , "000111100001001111111100011101" , "000111100001111111111100011100" , "000111100010101111111100011100" , "000111100011100111111100011011" , "000111100100010111111100011010" , "000111100101000111111100011001" , "000111100101110111111100011001"
, "000111100110101111111100011000" , "000111100111011111111100010111" , "000111101000001111111100010110" , "000111101000111111111100010110" , "000111101001110111111100010101" , "000111101010100111111100010100" , "000111101011010111111100010011" , "000111101100000111111100010011" , "000111101100111111111100010010" , "000111101101101111111100010001"
, "000111101110011111111100010000" , "000111101111001111111100010000" , "000111101111111111111100001111" , "000111110000110111111100001110" , "000111110001100111111100001101" , "000111110010010111111100001101" , "000111110011000111111100001100" , "000111110011111111111100001011" , "000111110100101111111100001010" , "000111110101011111111100001010"
, "000111110110001111111100001001" , "000111110111000111111100001000" , "000111110111110111111100000111" , "000111111000100111111100000110" , "000111111001010111111100000110" , "000111111010001111111100000101" , "000111111010111111111100000100" , "000111111011101111111100000011" , "000111111100011111111100000011" , "000111111101010111111100000010"
, "000111111110000111111100000001" , "000111111110110111111100000000" , "000111111111100111111011111111" , "001000000000010111111011111111" , "001000000001001111111011111110" , "001000000001111111111011111101" , "001000000010101111111011111100" , "001000000011011111111011111100" , "001000000100010111111011111011" , "001000000101000111111011111010"
, "001000000101110111111011111001" , "001000000110100111111011111000" , "001000000111011111111011111000" , "001000001000001111111011110111" , "001000001000111111111011110110" , "001000001001101111111011110101" , "001000001010011111111011110100" , "001000001011010111111011110100" , "001000001100000111111011110011" , "001000001100110111111011110010"
, "001000001101100111111011110001" , "001000001110011111111011110000" , "001000001111001111111011110000" , "001000001111111111111011101111" , "001000010000101111111011101110" , "001000010001100111111011101101" , "001000010010010111111011101100" , "001000010011000111111011101011" , "001000010011110111111011101011" , "001000010100100111111011101010"
, "001000010101011111111011101001" , "001000010110001111111011101000" , "001000010110111111111011100111" , "001000010111101111111011100111" , "001000011000100111111011100110" , "001000011001010111111011100101" , "001000011010000111111011100100" , "001000011010110111111011100011" , "001000011011101111111011100010" , "001000011100011111111011100010"
, "001000011101001111111011100001" , "001000011101111111111011100000" , "001000011110101111111011011111" , "001000011111100111111011011110" , "001000100000010111111011011101" , "001000100001000111111011011101" , "001000100001110111111011011100" , "001000100010101111111011011011" , "001000100011011111111011011010" , "001000100100001111111011011001"
, "001000100100111111111011011000" , "001000100101101111111011011000" , "001000100110100111111011010111" , "001000100111010111111011010110" , "001000101000000111111011010101" , "001000101000110111111011010100" , "001000101001101111111011010011" , "001000101010011111111011010011" , "001000101011001111111011010010" , "001000101011111111111011010001"
, "001000101100110111111011010000" , "001000101101100111111011001111" , "001000101110010111111011001110" , "001000101111000111111011001101" , "001000101111110111111011001101" , "001000110000101111111011001100" , "001000110001011111111011001011" , "001000110010001111111011001010" , "001000110010111111111011001001" , "001000110011110111111011001000"
, "001000110100100111111011000111" , "001000110101010111111011000110" , "001000110110000111111011000110" , "001000110110110111111011000101" , "001000110111101111111011000100" , "001000111000011111111011000011" , "001000111001001111111011000010" , "001000111001111111111011000001" , "001000111010110111111011000000" , "001000111011100111111011000000"
, "001000111100010111111010111111" , "001000111101000111111010111110" , "001000111101110111111010111101" , "001000111110101111111010111100" , "001000111111011111111010111011" , "001001000000001111111010111010" , "001001000000111111111010111001" , "001001000001110111111010111000" , "001001000010100111111010111000" , "001001000011010111111010110111"
, "001001000100000111111010110110" , "001001000100110111111010110101" , "001001000101101111111010110100" , "001001000110011111111010110011" , "001001000111001111111010110010" , "001001000111111111111010110001" , "001001001000110111111010110000" , "001001001001100111111010110000" , "001001001010010111111010101111" , "001001001011000111111010101110"
, "001001001011110111111010101101" , "001001001100101111111010101100" , "001001001101011111111010101011" , "001001001110001111111010101010" , "001001001110111111111010101001" , "001001001111101111111010101000" , "001001010000100111111010100111" , "001001010001010111111010100110" , "001001010010000111111010100110" , "001001010010110111111010100101"
, "001001010011101111111010100100" , "001001010100011111111010100011" , "001001010101001111111010100010" , "001001010101111111111010100001" , "001001010110101111111010100000" , "001001010111100111111010011111" , "001001011000010111111010011110" , "001001011001000111111010011101" , "001001011001110111111010011100" , "001001011010100111111010011011"
, "001001011011011111111010011011" , "001001011100001111111010011010" , "001001011100111111111010011001" , "001001011101101111111010011000" , "001001011110100111111010010111" , "001001011111010111111010010110" , "001001100000000111111010010101" , "001001100000110111111010010100" , "001001100001100111111010010011" , "001001100010011111111010010010"
, "001001100011001111111010010001" , "001001100011111111111010010000" , "001001100100101111111010001111" , "001001100101011111111010001110" , "001001100110010111111010001101" , "001001100111000111111010001101" , "001001100111110111111010001100" , "001001101000100111111010001011" , "001001101001011111111010001010" , "001001101010001111111010001001"
, "001001101010111111111010001000" , "001001101011101111111010000111" , "001001101100011111111010000110" , "001001101101010111111010000101" , "001001101110000111111010000100" , "001001101110110111111010000011" , "001001101111100111111010000010" , "001001110000010111111010000001" , "001001110001001111111010000000" , "001001110001111111111001111111"
, "001001110010101111111001111110" , "001001110011011111111001111101" , "001001110100001111111001111100" , "001001110101000111111001111011" , "001001110101110111111001111010" , "001001110110100111111001111001" , "001001110111010111111001111000" , "001001111000001111111001111000" , "001001111000111111111001110111" , "001001111001101111111001110110"
, "001001111010011111111001110101" , "001001111011001111111001110100" , "001001111100000111111001110011" , "001001111100110111111001110010" , "001001111101100111111001110001" , "001001111110010111111001110000" , "001001111111000111111001101111" , "001001111111111111111001101110" , "001010000000101111111001101101" , "001010000001011111111001101100"
, "001010000010001111111001101011" , "001010000010111111111001101010" , "001010000011110111111001101001" , "001010000100100111111001101000" , "001010000101010111111001100111" , "001010000110000111111001100110" , "001010000110110111111001100101" , "001010000111101111111001100100" , "001010001000011111111001100011" , "001010001001001111111001100010"
, "001010001001111111111001100001" , "001010001010101111111001100000" , "001010001011100111111001011111" , "001010001100010111111001011110" , "001010001101000111111001011101" , "001010001101110111111001011100" , "001010001110100111111001011011" , "001010001111011111111001011010" , "001010010000001111111001011001" , "001010010000111111111001011000"
, "001010010001101111111001010111" , "001010010010011111111001010110" , "001010010011010111111001010101" , "001010010100000111111001010100" , "001010010100110111111001010011" , "001010010101100111111001010010" , "001010010110010111111001010001" , "001010010111001111111001010000" , "001010010111111111111001001111" , "001010011000101111111001001110"
, "001010011001011111111001001101" , "001010011010001111111001001100" , "001010011011000111111001001011" , "001010011011110111111001001010" , "001010011100100111111001001001" , "001010011101010111111001001000" , "001010011110000111111001000111" , "001010011110111111111001000110" , "001010011111101111111001000101" , "001010100000011111111001000011"
, "001010100001001111111001000010" , "001010100001111111111001000001" , "001010100010110111111001000000" , "001010100011100111111000111111" , "001010100100010111111000111110" , "001010100101000111111000111101" , "001010100101110111111000111100" , "001010100110101111111000111011" , "001010100111011111111000111010" , "001010101000001111111000111001"
, "001010101000111111111000111000" , "001010101001101111111000110111" , "001010101010100111111000110110" , "001010101011010111111000110101" , "001010101100000111111000110100" , "001010101100110111111000110011" , "001010101101100111111000110010" , "001010101110011111111000110001" , "001010101111001111111000110000" , "001010101111111111111000101111"
, "001010110000101111111000101110" , "001010110001011111111000101101" , "001010110010010111111000101011" , "001010110011000111111000101010" , "001010110011110111111000101001" , "001010110100100111111000101000" , "001010110101010111111000100111" , "001010110110001111111000100110" , "001010110110111111111000100101" , "001010110111101111111000100100"
, "001010111000011111111000100011" , "001010111001001111111000100010" , "001010111010000111111000100001" , "001010111010110111111000100000" , "001010111011100111111000011111" , "001010111100010111111000011110" , "001010111101000111111000011101" , "001010111101110111111000011011" , "001010111110101111111000011010" , "001010111111011111111000011001"
, "001011000000001111111000011000" , "001011000000111111111000010111" , "001011000001101111111000010110" , "001011000010100111111000010101" , "001011000011010111111000010100" , "001011000100000111111000010011" , "001011000100110111111000010010" , "001011000101100111111000010001" , "001011000110011111111000010000" , "001011000111001111111000001110"
, "001011000111111111111000001101" , "001011001000101111111000001100" , "001011001001011111111000001011" , "001011001010001111111000001010" , "001011001011000111111000001001" , "001011001011110111111000001000" , "001011001100100111111000000111" , "001011001101010111111000000110" , "001011001110000111111000000101" , "001011001110111111111000000011"
, "001011001111101111111000000010" , "001011010000011111111000000001" , "001011010001001111111000000000" , "001011010001111111110111111111" , "001011010010110111110111111110" , "001011010011100111110111111101" , "001011010100010111110111111100" , "001011010101000111110111111011" , "001011010101110111110111111001" , "001011010110100111110111111000"
, "001011010111011111110111110111" , "001011011000001111110111110110" , "001011011000111111110111110101" , "001011011001101111110111110100" , "001011011010011111110111110011" , "001011011011010111110111110010" , "001011011100000111110111110001" , "001011011100110111110111101111" , "001011011101100111110111101110" , "001011011110010111110111101101"
, "001011011111000111110111101100" , "001011011111111111110111101011" , "001011100000101111110111101010" , "001011100001011111110111101001" , "001011100010001111110111101000" , "001011100010111111110111100110" , "001011100011110111110111100101" , "001011100100100111110111100100" , "001011100101010111110111100011" , "001011100110000111110111100010"
, "001011100110110111110111100001" , "001011100111100111110111100000" , "001011101000011111110111011110" , "001011101001001111110111011101" , "001011101001111111110111011100" , "001011101010101111110111011011" , "001011101011011111110111011010" , "001011101100001111110111011001" , "001011101101000111110111011000" , "001011101101110111110111010110"
, "001011101110100111110111010101" , "001011101111010111110111010100" , "001011110000000111110111010011" , "001011110000111111110111010010" , "001011110001101111110111010001" , "001011110010011111110111001111" , "001011110011001111110111001110" , "001011110011111111110111001101" , "001011110100101111110111001100" , "001011110101100111110111001011"
, "001011110110010111110111001010" , "001011110111000111110111001001" , "001011110111110111110111000111" , "001011111000100111110111000110" , "001011111001010111110111000101" , "001011111010001111110111000100" , "001011111010111111110111000011" , "001011111011101111110111000010" , "001011111100011111110111000000" , "001011111101001111110110111111"
, "001011111110000111110110111110" , "001011111110110111110110111101" , "001011111111100111110110111100" , "001100000000010111110110111010" , "001100000001000111110110111001" , "001100000001110111110110111000" , "001100000010101111110110110111" , "001100000011011111110110110110" , "001100000100001111110110110101" , "001100000100111111110110110011"
, "001100000101101111110110110010" , "001100000110011111110110110001" , "001100000111010111110110110000" , "001100001000000111110110101111" , "001100001000110111110110101101" , "001100001001100111110110101100" , "001100001010010111110110101011" , "001100001011000111110110101010" , "001100001011111111110110101001" , "001100001100101111110110100111"
, "001100001101011111110110100110" , "001100001110001111110110100101" , "001100001110111111110110100100" , "001100001111101111110110100011" , "001100010000100111110110100001" , "001100010001010111110110100000" , "001100010010000111110110011111" , "001100010010110111110110011110" , "001100010011100111110110011101" , "001100010100010111110110011011"
, "001100010101001111110110011010" , "001100010101111111110110011001" , "001100010110101111110110011000" , "001100010111011111110110010111" , "001100011000001111110110010101" , "001100011000111111110110010100" , "001100011001110111110110010011" , "001100011010100111110110010010" , "001100011011010111110110010000" , "001100011100000111110110001111"
, "001100011100110111110110001110" , "001100011101100111110110001101" , "001100011110011111110110001100" , "001100011111001111110110001010" , "001100011111111111110110001001" , "001100100000101111110110001000" , "001100100001011111110110000111" , "001100100010001111110110000101" , "001100100011000111110110000100" , "001100100011110111110110000011"
, "001100100100100111110110000010" , "001100100101010111110110000001" , "001100100110000111110101111111" , "001100100110110111110101111110" , "001100100111100111110101111101" , "001100101000011111110101111100" , "001100101001001111110101111010" , "001100101001111111110101111001" , "001100101010101111110101111000" , "001100101011011111110101110111"
, "001100101100001111110101110101" , "001100101101000111110101110100" , "001100101101110111110101110011" , "001100101110100111110101110010" , "001100101111010111110101110000" , "001100110000000111110101101111" , "001100110000110111110101101110" , "001100110001101111110101101101" , "001100110010011111110101101011" , "001100110011001111110101101010"
, "001100110011111111110101101001" , "001100110100101111110101101000" , "001100110101011111110101100110" , "001100110110001111110101100101" , "001100110111000111110101100100" , "001100110111110111110101100011" , "001100111000100111110101100001" , "001100111001010111110101100000" , "001100111010000111110101011111" , "001100111010110111110101011101"
, "001100111011101111110101011100" , "001100111100011111110101011011" , "001100111101001111110101011010" , "001100111101111111110101011000" , "001100111110101111110101010111" , "001100111111011111110101010110" , "001101000000001111110101010101" , "001101000001000111110101010011" , "001101000001110111110101010010" , "001101000010100111110101010001"
, "001101000011010111110101001111" , "001101000100000111110101001110" , "001101000100110111110101001101" , "001101000101101111110101001100" , "001101000110011111110101001010" , "001101000111001111110101001001" , "001101000111111111110101001000" , "001101001000101111110101000110" , "001101001001011111110101000101" , "001101001010001111110101000100"
, "001101001011000111110101000011" , "001101001011110111110101000001" , "001101001100100111110101000000" , "001101001101010111110100111111" , "001101001110000111110100111101" , "001101001110110111110100111100" , "001101001111100111110100111011" , "001101010000011111110100111010" , "001101010001001111110100111000" , "001101010001111111110100110111"
, "001101010010101111110100110110" , "001101010011011111110100110100" , "001101010100001111110100110011" , "001101010101000111110100110010" , "001101010101110111110100110000" , "001101010110100111110100101111" , "001101010111010111110100101110" , "001101011000000111110100101100" , "001101011000110111110100101011" , "001101011001100111110100101010"
, "001101011010011111110100101000" , "001101011011001111110100100111" , "001101011011111111110100100110" , "001101011100101111110100100101" , "001101011101011111110100100011" , "001101011110001111110100100010" , "001101011110111111110100100001" , "001101011111110111110100011111" , "001101100000100111110100011110" , "001101100001010111110100011101"
, "001101100010000111110100011011" , "001101100010110111110100011010" , "001101100011100111110100011001" , "001101100100010111110100010111" , "001101100101001111110100010110" , "001101100101111111110100010101" , "001101100110101111110100010011" , "001101100111011111110100010010" , "001101101000001111110100010001" , "001101101000111111110100001111"
, "001101101001101111110100001110" , "001101101010011111110100001101" , "001101101011010111110100001011" , "001101101100000111110100001010" , "001101101100110111110100001001" , "001101101101100111110100000111" , "001101101110010111110100000110" , "001101101111000111110100000101" , "001101101111110111110100000011" , "001101110000101111110100000010"
, "001101110001011111110100000000" , "001101110010001111110011111111" , "001101110010111111110011111110" , "001101110011101111110011111100" , "001101110100011111110011111011" , "001101110101001111110011111010" , "001101110110000111110011111000" , "001101110110110111110011110111" , "001101110111100111110011110110" , "001101111000010111110011110100"
, "001101111001000111110011110011" , "001101111001110111110011110010" , "001101111010100111110011110000" , "001101111011010111110011101111" , "001101111100001111110011101101" , "001101111100111111110011101100" , "001101111101101111110011101011" , "001101111110011111110011101001" , "001101111111001111110011101000" , "001101111111111111110011100111"
, "001110000000101111110011100101" , "001110000001100111110011100100" , "001110000010010111110011100010" , "001110000011000111110011100001" , "001110000011110111110011100000" , "001110000100100111110011011110" , "001110000101010111110011011101" , "001110000110000111110011011100" , "001110000110110111110011011010" , "001110000111101111110011011001"
, "001110001000011111110011010111" , "001110001001001111110011010110" , "001110001001111111110011010101" , "001110001010101111110011010011" , "001110001011011111110011010010" , "001110001100001111110011010000" , "001110001100111111110011001111" , "001110001101110111110011001110" , "001110001110100111110011001100" , "001110001111010111110011001011"
, "001110010000000111110011001001" , "001110010000110111110011001000" , "001110010001100111110011000111" , "001110010010010111110011000101" , "001110010011000111110011000100" , "001110010011111111110011000010" , "001110010100101111110011000001" , "001110010101011111110011000000" , "001110010110001111110010111110" , "001110010110111111110010111101"
, "001110010111101111110010111011" , "001110011000011111110010111010" , "001110011001001111110010111001" , "001110011010000111110010110111" , "001110011010110111110010110110" , "001110011011100111110010110100" , "001110011100010111110010110011" , "001110011101000111110010110001" , "001110011101110111110010110000" , "001110011110100111110010101111"
, "001110011111010111110010101101" , "001110100000001111110010101100" , "001110100000111111110010101010" , "001110100001101111110010101001" , "001110100010011111110010101000" , "001110100011001111110010100110" , "001110100011111111110010100101" , "001110100100101111110010100011" , "001110100101011111110010100010" , "001110100110001111110010100000"
, "001110100111000111110010011111" , "001110100111110111110010011110" , "001110101000100111110010011100" , "001110101001010111110010011011" , "001110101010000111110010011001" , "001110101010110111110010011000" , "001110101011100111110010010110" , "001110101100010111110010010101" , "001110101101001111110010010011" , "001110101101111111110010010010"
, "001110101110101111110010010001" , "001110101111011111110010001111" , "001110110000001111110010001110" , "001110110000111111110010001100" , "001110110001101111110010001011" , "001110110010011111110010001001" , "001110110011001111110010001000" , "001110110100000111110010000110" , "001110110100110111110010000101" , "001110110101100111110010000011"
, "001110110110010111110010000010" , "001110110111000111110010000001" , "001110110111110111110001111111" , "001110111000100111110001111110" , "001110111001010111110001111100" , "001110111010000111110001111011" , "001110111010111111110001111001" , "001110111011101111110001111000" , "001110111100011111110001110110" , "001110111101001111110001110101"
, "001110111101111111110001110011" , "001110111110101111110001110010" , "001110111111011111110001110000" , "001111000000001111110001101111" , "001111000000111111110001101110" , "001111000001110111110001101100" , "001111000010100111110001101011" , "001111000011010111110001101001" , "001111000100000111110001101000" , "001111000100110111110001100110"
, "001111000101100111110001100101" , "001111000110010111110001100011" , "001111000111000111110001100010" , "001111000111110111110001100000" , "001111001000100111110001011111" , "001111001001011111110001011101" , "001111001010001111110001011100" , "001111001010111111110001011010" , "001111001011101111110001011001" , "001111001100011111110001010111"
, "001111001101001111110001010110" , "001111001101111111110001010100" , "001111001110101111110001010011" , "001111001111011111110001010001" , "001111010000010111110001010000" , "001111010001000111110001001110" , "001111010001110111110001001101" , "001111010010100111110001001011" , "001111010011010111110001001010" , "001111010100000111110001001000"
, "001111010100110111110001000111" , "001111010101100111110001000101" , "001111010110010111110001000100" , "001111010111000111110001000010" , "001111010111111111110001000001" , "001111011000101111110000111111" , "001111011001011111110000111110" , "001111011010001111110000111100" , "001111011010111111110000111011" , "001111011011101111110000111001"
, "001111011100011111110000111000" , "001111011101001111110000110110" , "001111011101111111110000110101" , "001111011110101111110000110011" , "001111011111011111110000110010" , "001111100000010111110000110000" , "001111100001000111110000101111" , "001111100001110111110000101101" , "001111100010100111110000101100" , "001111100011010111110000101010"
, "001111100100000111110000101000" , "001111100100110111110000100111" , "001111100101100111110000100101" , "001111100110010111110000100100" , "001111100111000111110000100010" , "001111100111111111110000100001" , "001111101000101111110000011111" , "001111101001011111110000011110" , "001111101010001111110000011100" , "001111101010111111110000011011"
, "001111101011101111110000011001" , "001111101100011111110000011000" , "001111101101001111110000010110" , "001111101101111111110000010100" , "001111101110101111110000010011" , "001111101111011111110000010001" , "001111110000010111110000010000" , "001111110001000111110000001110" , "001111110001110111110000001101" , "001111110010100111110000001011"
, "001111110011010111110000001010" , "001111110100000111110000001000" , "001111110100110111110000000111" , "001111110101100111110000000101" , "001111110110010111110000000011" , "001111110111000111110000000010" , "001111110111110111110000000000" , "001111111000101111101111111111" , "001111111001011111101111111101" , "001111111010001111101111111100"
, "001111111010111111101111111010" , "001111111011101111101111111001" , "001111111100011111101111110111" , "001111111101001111101111110101" , "001111111101111111101111110100" , "001111111110101111101111110010" , "001111111111011111101111110001" , "010000000000001111101111101111" , "010000000000111111101111101110" , "010000000001110111101111101100"
, "010000000010100111101111101010" , "010000000011010111101111101001" , "010000000100000111101111100111" , "010000000100110111101111100110" , "010000000101100111101111100100" , "010000000110010111101111100011" , "010000000111000111101111100001" , "010000000111110111101111011111" , "010000001000100111101111011110" , "010000001001010111101111011100"
, "010000001010000111101111011011" , "010000001010111111101111011001" , "010000001011101111101111010111" , "010000001100011111101111010110" , "010000001101001111101111010100" , "010000001101111111101111010011" , "010000001110101111101111010001" , "010000001111011111101111001111" , "010000010000001111101111001110" , "010000010000111111101111001100"
, "010000010001101111101111001011" , "010000010010011111101111001001" , "010000010011001111101111000111" , "010000010011111111101111000110" , "010000010100110111101111000100" , "010000010101100111101111000011" , "010000010110010111101111000001" , "010000010111000111101110111111" , "010000010111110111101110111110" , "010000011000100111101110111100"
, "010000011001010111101110111011" , "010000011010000111101110111001" , "010000011010110111101110110111" , "010000011011100111101110110110" , "010000011100010111101110110100" , "010000011101000111101110110011" , "010000011101110111101110110001" , "010000011110100111101110101111" , "010000011111011111101110101110" , "010000100000001111101110101100"
, "010000100000111111101110101010" , "010000100001101111101110101001" , "010000100010011111101110100111" , "010000100011001111101110100110" , "010000100011111111101110100100" , "010000100100101111101110100010" , "010000100101011111101110100001" , "010000100110001111101110011111" , "010000100110111111101110011101" , "010000100111101111101110011100"
, "010000101000011111101110011010" , "010000101001001111101110011001" , "010000101010000111101110010111" , "010000101010110111101110010101" , "010000101011100111101110010100" , "010000101100010111101110010010" , "010000101101000111101110010000" , "010000101101110111101110001111" , "010000101110100111101110001101" , "010000101111010111101110001011"
, "010000110000000111101110001010" , "010000110000110111101110001000" , "010000110001100111101110000111" , "010000110010010111101110000101" , "010000110011000111101110000011" , "010000110011110111101110000010" , "010000110100100111101110000000" , "010000110101010111101101111110" , "010000110110001111101101111101" , "010000110110111111101101111011"
, "010000110111101111101101111001" , "010000111000011111101101111000" , "010000111001001111101101110110" , "010000111001111111101101110100" , "010000111010101111101101110011" , "010000111011011111101101110001" , "010000111100001111101101101111" , "010000111100111111101101101110" , "010000111101101111101101101100" , "010000111110011111101101101010"
, "010000111111001111101101101001" , "010000111111111111101101100111" , "010001000000101111101101100101" , "010001000001011111101101100100" , "010001000010001111101101100010" , "010001000011000111101101100000" , "010001000011110111101101011111" , "010001000100100111101101011101" , "010001000101010111101101011011" , "010001000110000111101101011010"
, "010001000110110111101101011000" , "010001000111100111101101010110" , "010001001000010111101101010101" , "010001001001000111101101010011" , "010001001001110111101101010001" , "010001001010100111101101010000" , "010001001011010111101101001110" , "010001001100000111101101001100" , "010001001100110111101101001011" , "010001001101100111101101001001"
, "010001001110010111101101000111" , "010001001111000111101101000101" , "010001001111110111101101000100" , "010001010000100111101101000010" , "010001010001011111101101000000" , "010001010010001111101100111111" , "010001010010111111101100111101" , "010001010011101111101100111011" , "010001010100011111101100111010" , "010001010101001111101100111000"
, "010001010101111111101100110110" , "010001010110101111101100110100" , "010001010111011111101100110011" , "010001011000001111101100110001" , "010001011000111111101100101111" , "010001011001101111101100101110" , "010001011010011111101100101100" , "010001011011001111101100101010" , "010001011011111111101100101001" , "010001011100101111101100100111"
, "010001011101011111101100100101" , "010001011110001111101100100011" , "010001011110111111101100100010" , "010001011111101111101100100000" , "010001100000011111101100011110" , "010001100001010111101100011100" , "010001100010000111101100011011" , "010001100010110111101100011001" , "010001100011100111101100010111" , "010001100100010111101100010110"
, "010001100101000111101100010100" , "010001100101110111101100010010" , "010001100110100111101100010000" , "010001100111010111101100001111" , "010001101000000111101100001101" , "010001101000110111101100001011" , "010001101001100111101100001010" , "010001101010010111101100001000" , "010001101011000111101100000110" , "010001101011110111101100000100"
, "010001101100100111101100000011" , "010001101101010111101100000001" , "010001101110000111101011111111" , "010001101110110111101011111101" , "010001101111100111101011111100" , "010001110000010111101011111010" , "010001110001000111101011111000" , "010001110001110111101011110110" , "010001110010100111101011110101" , "010001110011010111101011110011"
, "010001110100000111101011110001" , "010001110100111111101011101111" , "010001110101101111101011101110" , "010001110110011111101011101100" , "010001110111001111101011101010" , "010001110111111111101011101000" , "010001111000101111101011100111" , "010001111001011111101011100101" , "010001111010001111101011100011" , "010001111010111111101011100001"
, "010001111011101111101011100000" , "010001111100011111101011011110" , "010001111101001111101011011100" , "010001111101111111101011011010" , "010001111110101111101011011001" , "010001111111011111101011010111" , "010010000000001111101011010101" , "010010000000111111101011010011" , "010010000001101111101011010001" , "010010000010011111101011010000"
, "010010000011001111101011001110" , "010010000011111111101011001100" , "010010000100101111101011001010" , "010010000101011111101011001001" , "010010000110001111101011000111" , "010010000110111111101011000101" , "010010000111101111101011000011" , "010010001000011111101011000001" , "010010001001001111101011000000" , "010010001001111111101010111110"
, "010010001010101111101010111100" , "010010001011011111101010111010" , "010010001100001111101010111001" , "010010001100111111101010110111" , "010010001101101111101010110101" , "010010001110100111101010110011" , "010010001111010111101010110001" , "010010010000000111101010110000" , "010010010000110111101010101110" , "010010010001100111101010101100"
, "010010010010010111101010101010" , "010010010011000111101010101000" , "010010010011110111101010100111" , "010010010100100111101010100101" , "010010010101010111101010100011" , "010010010110000111101010100001" , "010010010110110111101010011111" , "010010010111100111101010011110" , "010010011000010111101010011100" , "010010011001000111101010011010"
, "010010011001110111101010011000" , "010010011010100111101010010110" , "010010011011010111101010010101" , "010010011100000111101010010011" , "010010011100110111101010010001" , "010010011101100111101010001111" , "010010011110010111101010001101" , "010010011111000111101010001100" , "010010011111110111101010001010" , "010010100000100111101010001000"
, "010010100001010111101010000110" , "010010100010000111101010000100" , "010010100010110111101010000010" , "010010100011100111101010000001" , "010010100100010111101001111111" , "010010100101000111101001111101" , "010010100101110111101001111011" , "010010100110100111101001111001" , "010010100111010111101001111000" , "010010101000000111101001110110"
, "010010101000110111101001110100" , "010010101001100111101001110010" , "010010101010010111101001110000" , "010010101011000111101001101110" , "010010101011110111101001101101" , "010010101100100111101001101011" , "010010101101010111101001101001" , "010010101110000111101001100111" , "010010101110110111101001100101" , "010010101111100111101001100011"
, "010010110000010111101001100010" , "010010110001000111101001100000" , "010010110001110111101001011110" , "010010110010100111101001011100" , "010010110011010111101001011010" , "010010110100000111101001011000" , "010010110100110111101001010110" , "010010110101100111101001010101" , "010010110110010111101001010011" , "010010110111000111101001010001"
, "010010110111110111101001001111" , "010010111000100111101001001101" , "010010111001010111101001001011" , "010010111010000111101001001001" , "010010111010110111101001001000" , "010010111011100111101001000110" , "010010111100010111101001000100" , "010010111101000111101001000010" , "010010111101110111101001000000" , "010010111110100111101000111110"
, "010010111111010111101000111100" , "010011000000000111101000111011" , "010011000000110111101000111001" , "010011000001100111101000110111" , "010011000010010111101000110101" , "010011000011000111101000110011" , "010011000011110111101000110001" , "010011000100100111101000101111" , "010011000101010111101000101110" , "010011000110000111101000101100"
, "010011000110110111101000101010" , "010011000111100111101000101000" , "010011001000010111101000100110" , "010011001001000111101000100100" , "010011001001110111101000100010" , "010011001010100111101000100000" , "010011001011010111101000011111" , "010011001100000111101000011101" , "010011001100110111101000011011" , "010011001101100111101000011001"
, "010011001110010111101000010111" , "010011001111000111101000010101" , "010011001111110111101000010011" , "010011010000100111101000010001" , "010011010001010111101000001111" , "010011010010000111101000001110" , "010011010010110111101000001100" , "010011010011100111101000001010" , "010011010100010111101000001000" , "010011010101000111101000000110"
, "010011010101110111101000000100" , "010011010110100111101000000010" , "010011010111010111101000000000" , "010011011000000111100111111110" , "010011011000110111100111111100" , "010011011001100111100111111011" , "010011011010010111100111111001" , "010011011011000111100111110111" , "010011011011110111100111110101" , "010011011100100111100111110011"
, "010011011101010111100111110001" , "010011011110000111100111101111" , "010011011110110111100111101101" , "010011011111100111100111101011" , "010011100000010111100111101001" , "010011100001000111100111100111" , "010011100001110111100111100110" , "010011100010100111100111100100" , "010011100011010111100111100010" , "010011100100000111100111100000"
, "010011100100110111100111011110" , "010011100101100111100111011100" , "010011100110010111100111011010" , "010011100111000111100111011000" , "010011100111110111100111010110" , "010011101000100111100111010100" , "010011101001010111100111010010" , "010011101010000111100111010000" , "010011101010110111100111001110" , "010011101011100111100111001100"
, "010011101100010111100111001011" , "010011101101000111100111001001" , "010011101101110111100111000111" , "010011101110100111100111000101" , "010011101111010111100111000011" , "010011110000000111100111000001" , "010011110000110111100110111111" , "010011110001011111100110111101" , "010011110010001111100110111011" , "010011110010111111100110111001"
, "010011110011101111100110110111" , "010011110100011111100110110101" , "010011110101001111100110110011" , "010011110101111111100110110001" , "010011110110101111100110101111" , "010011110111011111100110101101" , "010011111000001111100110101011" , "010011111000111111100110101010" , "010011111001101111100110101000" , "010011111010011111100110100110"
, "010011111011001111100110100100" , "010011111011111111100110100010" , "010011111100101111100110100000" , "010011111101011111100110011110" , "010011111110001111100110011100" , "010011111110111111100110011010" , "010011111111101111100110011000" , "010100000000011111100110010110" , "010100000001001111100110010100" , "010100000001111111100110010010"
, "010100000010101111100110010000" , "010100000011011111100110001110" , "010100000100001111100110001100" , "010100000100111111100110001010" , "010100000101101111100110001000" , "010100000110011111100110000110" , "010100000111001111100110000100" , "010100000111111111100110000010" , "010100001000101111100110000000" , "010100001001011111100101111110"
, "010100001010000111100101111100" , "010100001010110111100101111010" , "010100001011100111100101111000" , "010100001100010111100101110110" , "010100001101000111100101110100" , "010100001101110111100101110010" , "010100001110100111100101110000" , "010100001111010111100101101110" , "010100010000000111100101101100" , "010100010000110111100101101010"
, "010100010001100111100101101000" , "010100010010010111100101100110" , "010100010011000111100101100100" , "010100010011110111100101100010" , "010100010100100111100101100000" , "010100010101010111100101011111" , "010100010110000111100101011101" , "010100010110110111100101011011" , "010100010111100111100101011001" , "010100011000010111100101010111"
, "010100011001000111100101010101" , "010100011001110111100101010011" , "010100011010100111100101010001" , "010100011011010111100101001110" , "010100011011111111100101001100" , "010100011100101111100101001010" , "010100011101011111100101001000" , "010100011110001111100101000110" , "010100011110111111100101000100" , "010100011111101111100101000010"
, "010100100000011111100101000000" , "010100100001001111100100111110" , "010100100001111111100100111100" , "010100100010101111100100111010" , "010100100011011111100100111000" , "010100100100001111100100110110" , "010100100100111111100100110100" , "010100100101101111100100110010" , "010100100110011111100100110000" , "010100100111001111100100101110"
, "010100100111111111100100101100" , "010100101000101111100100101010" , "010100101001011111100100101000" , "010100101010001111100100100110" , "010100101010110111100100100100" , "010100101011100111100100100010" , "010100101100010111100100100000" , "010100101101000111100100011110" , "010100101101110111100100011100" , "010100101110100111100100011010"
, "010100101111010111100100011000" , "010100110000000111100100010110" , "010100110000110111100100010100" , "010100110001100111100100010010" , "010100110010010111100100010000" , "010100110011000111100100001110" , "010100110011110111100100001100" , "010100110100100111100100001010" , "010100110101010111100100001000" , "010100110110000111100100000110"
, "010100110110110111100100000100" , "010100110111100111100100000001" , "010100111000001111100011111111" , "010100111000111111100011111101" , "010100111001101111100011111011" , "010100111010011111100011111001" , "010100111011001111100011110111" , "010100111011111111100011110101" , "010100111100101111100011110011" , "010100111101011111100011110001"
, "010100111110001111100011101111" , "010100111110111111100011101101" , "010100111111101111100011101011" , "010101000000011111100011101001" , "010101000001001111100011100111" , "010101000001111111100011100101" , "010101000010101111100011100011" , "010101000011011111100011100001" , "010101000100000111100011011110" , "010101000100110111100011011100"
, "010101000101100111100011011010" , "010101000110010111100011011000" , "010101000111000111100011010110" , "010101000111110111100011010100" , "010101001000100111100011010010" , "010101001001010111100011010000" , "010101001010000111100011001110" , "010101001010110111100011001100" , "010101001011100111100011001010" , "010101001100010111100011001000"
, "010101001101000111100011000110" , "010101001101110111100011000100" , "010101001110011111100011000001" , "010101001111001111100010111111" , "010101001111111111100010111101" , "010101010000101111100010111011" , "010101010001011111100010111001" , "010101010010001111100010110111" , "010101010010111111100010110101" , "010101010011101111100010110011"
, "010101010100011111100010110001" , "010101010101001111100010101111" , "010101010101111111100010101101" , "010101010110101111100010101010" , "010101010111011111100010101000" , "010101011000001111100010100110" , "010101011000110111100010100100" , "010101011001100111100010100010" , "010101011010010111100010100000" , "010101011011000111100010011110"
, "010101011011110111100010011100" , "010101011100100111100010011010" , "010101011101010111100010011000" , "010101011110000111100010010101" , "010101011110110111100010010011" , "010101011111100111100010010001" , "010101100000010111100010001111" , "010101100001000111100010001101" , "010101100001101111100010001011" , "010101100010011111100010001001"
, "010101100011001111100010000111" , "010101100011111111100010000101" , "010101100100101111100010000010" , "010101100101011111100010000000" , "010101100110001111100001111110" , "010101100110111111100001111100" , "010101100111101111100001111010" , "010101101000011111100001111000" , "010101101001001111100001110110" , "010101101001111111100001110100"
, "010101101010100111100001110001" , "010101101011010111100001101111" , "010101101100000111100001101101" , "010101101100110111100001101011" , "010101101101100111100001101001" , "010101101110010111100001100111" , "010101101111000111100001100101" , "010101101111110111100001100011" , "010101110000100111100001100000" , "010101110001010111100001011110"
, "010101110010000111100001011100" , "010101110010101111100001011010" , "010101110011011111100001011000" , "010101110100001111100001010110" , "010101110100111111100001010100" , "010101110101101111100001010001" , "010101110110011111100001001111" , "010101110111001111100001001101" , "010101110111111111100001001011" , "010101111000101111100001001001"
, "010101111001011111100001000111" , "010101111010000111100001000101" , "010101111010110111100001000010" , "010101111011100111100001000000" , "010101111100010111100000111110" , "010101111101000111100000111100" , "010101111101110111100000111010" , "010101111110100111100000111000" , "010101111111010111100000110101" , "010110000000000111100000110011"
, "010110000000110111100000110001" , "010110000001100111100000101111" , "010110000010001111100000101101" , "010110000010111111100000101011" , "010110000011101111100000101000" , "010110000100011111100000100110" , "010110000101001111100000100100" , "010110000101111111100000100010" , "010110000110101111100000100000" , "010110000111011111100000011110"
, "010110001000001111100000011011" , "010110001000110111100000011001" , "010110001001100111100000010111" , "010110001010010111100000010101" , "010110001011000111100000010011" , "010110001011110111100000010001" , "010110001100100111100000001110" , "010110001101010111100000001100" , "010110001110000111100000001010" , "010110001110110111100000001000"
, "010110001111100111100000000110" , "010110010000001111100000000011" , "010110010000111111100000000001" , "010110010001101111011111111111" , "010110010010011111011111111101" , "010110010011001111011111111011" , "010110010011111111011111111001" , "010110010100101111011111110110" , "010110010101011111011111110100" , "010110010110001111011111110010"
, "010110010110110111011111110000" , "010110010111100111011111101110" , "010110011000010111011111101011" , "010110011001000111011111101001" , "010110011001110111011111100111" , "010110011010100111011111100101" , "010110011011010111011111100011" , "010110011100000111011111100000" , "010110011100110111011111011110" , "010110011101011111011111011100"
, "010110011110001111011111011010" , "010110011110111111011111011000" , "010110011111101111011111010101" , "010110100000011111011111010011" , "010110100001001111011111010001" , "010110100001111111011111001111" , "010110100010101111011111001101" , "010110100011010111011111001010" , "010110100100000111011111001000" , "010110100100110111011111000110"
, "010110100101100111011111000100" , "010110100110010111011111000001" , "010110100111000111011110111111" , "010110100111110111011110111101" , "010110101000100111011110111011" , "010110101001001111011110111001" , "010110101001111111011110110110" , "010110101010101111011110110100" , "010110101011011111011110110010" , "010110101100001111011110110000"
, "010110101100111111011110101101" , "010110101101101111011110101011" , "010110101110011111011110101001" , "010110101111000111011110100111" , "010110101111110111011110100100" , "010110110000100111011110100010" , "010110110001010111011110100000" , "010110110010000111011110011110" , "010110110010110111011110011100" , "010110110011100111011110011001"
, "010110110100010111011110010111" , "010110110100111111011110010101" , "010110110101101111011110010011" , "010110110110011111011110010000" , "010110110111001111011110001110" , "010110110111111111011110001100" , "010110111000101111011110001010" , "010110111001011111011110000111" , "010110111010001111011110000101" , "010110111010110111011110000011"
, "010110111011100111011110000001" , "010110111100010111011101111110" , "010110111101000111011101111100" , "010110111101110111011101111010" , "010110111110100111011101111000" , "010110111111010111011101110101" , "010110111111111111011101110011" , "010111000000101111011101110001" , "010111000001011111011101101111" , "010111000010001111011101101100"
, "010111000010111111011101101010" , "010111000011101111011101101000" , "010111000100011111011101100110" , "010111000101000111011101100011" , "010111000101110111011101100001" , "010111000110100111011101011111" , "010111000111010111011101011100" , "010111001000000111011101011010" , "010111001000110111011101011000" , "010111001001100111011101010110"
, "010111001010001111011101010011" , "010111001010111111011101010001" , "010111001011101111011101001111" , "010111001100011111011101001101" , "010111001101001111011101001010" , "010111001101111111011101001000" , "010111001110101111011101000110" , "010111001111010111011101000011" , "010111010000000111011101000001" , "010111010000110111011100111111"
, "010111010001100111011100111101" , "010111010010010111011100111010" , "010111010011000111011100111000" , "010111010011110111011100110110" , "010111010100011111011100110011" , "010111010101001111011100110001" , "010111010101111111011100101111" , "010111010110101111011100101101" , "010111010111011111011100101010" , "010111011000001111011100101000"
, "010111011000111111011100100110" , "010111011001100111011100100011" , "010111011010010111011100100001" , "010111011011000111011100011111" , "010111011011110111011100011100" , "010111011100100111011100011010" , "010111011101010111011100011000" , "010111011101111111011100010110" , "010111011110101111011100010011" , "010111011111011111011100010001"
, "010111100000001111011100001111" , "010111100000111111011100001100" , "010111100001101111011100001010" , "010111100010011111011100001000" , "010111100011000111011100000101" , "010111100011110111011100000011" , "010111100100100111011100000001" , "010111100101010111011011111110" , "010111100110000111011011111100" , "010111100110110111011011111010"
, "010111100111011111011011111000" , "010111101000001111011011110101" , "010111101000111111011011110011" , "010111101001101111011011110001" , "010111101010011111011011101110" , "010111101011001111011011101100" , "010111101011110111011011101010" , "010111101100100111011011100111" , "010111101101010111011011100101" , "010111101110000111011011100011"
, "010111101110110111011011100000" , "010111101111100111011011011110" , "010111110000001111011011011100" , "010111110000111111011011011001" , "010111110001101111011011010111" , "010111110010011111011011010101" , "010111110011001111011011010010" , "010111110011111111011011010000" , "010111110100100111011011001110" , "010111110101010111011011001011"
, "010111110110000111011011001001" , "010111110110110111011011000111" , "010111110111100111011011000100" , "010111111000010111011011000010" , "010111111000111111011011000000" , "010111111001101111011010111101" , "010111111010011111011010111011" , "010111111011001111011010111001" , "010111111011111111011010110110" , "010111111100101111011010110100"
, "010111111101010111011010110001" , "010111111110000111011010101111" , "010111111110110111011010101101" , "010111111111100111011010101010" , "011000000000010111011010101000" , "011000000001000111011010100110" , "011000000001101111011010100011" , "011000000010011111011010100001" , "011000000011001111011010011111" , "011000000011111111011010011100"
, "011000000100101111011010011010" , "011000000101010111011010011000" , "011000000110000111011010010101" , "011000000110110111011010010011" , "011000000111100111011010010000" , "011000001000010111011010001110" , "011000001001000111011010001100" , "011000001001101111011010001001" , "011000001010011111011010000111" , "011000001011001111011010000101"
, "011000001011111111011010000010" , "011000001100101111011010000000" , "011000001101011111011001111101" , "011000001110000111011001111011" , "011000001110110111011001111001" , "011000001111100111011001110110" , "011000010000010111011001110100" , "011000010001000111011001110010" , "011000010001101111011001101111" , "011000010010011111011001101101"
, "011000010011001111011001101010" , "011000010011111111011001101000" , "011000010100101111011001100110" , "011000010101010111011001100011" , "011000010110000111011001100001" , "011000010110110111011001011110" , "011000010111100111011001011100" , "011000011000010111011001011010" , "011000011001000111011001010111" , "011000011001101111011001010101"
, "011000011010011111011001010010" , "011000011011001111011001010000" , "011000011011111111011001001110" , "011000011100101111011001001011" , "011000011101010111011001001001" , "011000011110000111011001000110" , "011000011110110111011001000100" , "011000011111100111011001000010" , "011000100000010111011000111111" , "011000100000111111011000111101"
, "011000100001101111011000111010" , "011000100010011111011000111000" , "011000100011001111011000110110" , "011000100011111111011000110011" , "011000100100100111011000110001" , "011000100101010111011000101110" , "011000100110000111011000101100" , "011000100110110111011000101010" , "011000100111100111011000100111" , "011000101000001111011000100101"
, "011000101000111111011000100010" , "011000101001101111011000100000" , "011000101010011111011000011101" , "011000101011001111011000011011" , "011000101011110111011000011001" , "011000101100100111011000010110" , "011000101101010111011000010100" , "011000101110000111011000010001" , "011000101110110111011000001111" , "011000101111011111011000001101"
, "011000110000001111011000001010" , "011000110000111111011000001000" , "011000110001101111011000000101" , "011000110010011111011000000011" , "011000110011000111011000000000" , "011000110011110111010111111110" , "011000110100100111010111111011" , "011000110101010111010111111001" , "011000110110000111010111110111" , "011000110110101111010111110100"
, "011000110111011111010111110010" , "011000111000001111010111101111" , "011000111000111111010111101101" , "011000111001100111010111101010" , "011000111010010111010111101000" , "011000111011000111010111100110" , "011000111011110111010111100011" , "011000111100100111010111100001" , "011000111101001111010111011110" , "011000111101111111010111011100"
, "011000111110101111010111011001" , "011000111111011111010111010111" , "011001000000001111010111010100" , "011001000000110111010111010010" , "011001000001100111010111001111" , "011001000010010111010111001101" , "011001000011000111010111001011" , "011001000011101111010111001000" , "011001000100011111010111000110" , "011001000101001111010111000011"
, "011001000101111111010111000001" , "011001000110101111010110111110" , "011001000111010111010110111100" , "011001001000000111010110111001" , "011001001000110111010110110111" , "011001001001100111010110110100" , "011001001010001111010110110010" , "011001001010111111010110101111" , "011001001011101111010110101101" , "011001001100011111010110101010"
, "011001001101001111010110101000" , "011001001101110111010110100110" , "011001001110100111010110100011" , "011001001111010111010110100001" , "011001010000000111010110011110" , "011001010000101111010110011100" , "011001010001011111010110011001" , "011001010010001111010110010111" , "011001010010111111010110010100" , "011001010011101111010110010010"
, "011001010100010111010110001111" , "011001010101000111010110001101" , "011001010101110111010110001010" , "011001010110100111010110001000" , "011001010111001111010110000101" , "011001010111111111010110000011" , "011001011000101111010110000000" , "011001011001011111010101111110" , "011001011010000111010101111011" , "011001011010110111010101111001"
, "011001011011100111010101110110" , "011001011100010111010101110100" , "011001011101000111010101110001" , "011001011101101111010101101111" , "011001011110011111010101101100" , "011001011111001111010101101010" , "011001011111111111010101100111" , "011001100000100111010101100101" , "011001100001010111010101100010" , "011001100010000111010101100000"
, "011001100010110111010101011101" , "011001100011011111010101011011" , "011001100100001111010101011000" , "011001100100111111010101010110" , "011001100101101111010101010011" , "011001100110010111010101010001" , "011001100111000111010101001110" , "011001100111110111010101001100" , "011001101000100111010101001001" , "011001101001001111010101000111"
, "011001101001111111010101000100" , "011001101010101111010101000010" , "011001101011011111010100111111" , "011001101100000111010100111101" , "011001101100110111010100111010" , "011001101101100111010100111000" , "011001101110010111010100110101" , "011001101110111111010100110010" , "011001101111101111010100110000" , "011001110000011111010100101101"
, "011001110001001111010100101011" , "011001110001110111010100101000" , "011001110010100111010100100110" , "011001110011010111010100100011" , "011001110100000111010100100001" , "011001110100101111010100011110" , "011001110101011111010100011100" , "011001110110001111010100011001" , "011001110110111111010100010111" , "011001110111100111010100010100"
, "011001111000010111010100010010" , "011001111001000111010100001111" , "011001111001110111010100001100" , "011001111010011111010100001010" , "011001111011001111010100000111" , "011001111011111111010100000101" , "011001111100101111010100000010" , "011001111101010111010100000000" , "011001111110000111010011111101" , "011001111110110111010011111011"
, "011001111111100111010011111000" , "011010000000001111010011110110" , "011010000000111111010011110011" , "011010000001101111010011110000" , "011010000010011111010011101110" , "011010000011000111010011101011" , "011010000011110111010011101001" , "011010000100100111010011100110" , "011010000101010111010011100100" , "011010000101111111010011100001"
, "011010000110101111010011011111" , "011010000111011111010011011100" , "011010001000001111010011011001" , "011010001000110111010011010111" , "011010001001100111010011010100" , "011010001010010111010011010010" , "011010001010111111010011001111" , "011010001011101111010011001101" , "011010001100011111010011001010" , "011010001101001111010011000111"
, "011010001101110111010011000101" , "011010001110100111010011000010" , "011010001111010111010011000000" , "011010010000000111010010111101" , "011010010000101111010010111011" , "011010010001011111010010111000" , "011010010010001111010010110101" , "011010010010111111010010110011" , "011010010011100111010010110000" , "011010010100010111010010101110"
, "011010010101000111010010101011" , "011010010101101111010010101000" , "011010010110011111010010100110" , "011010010111001111010010100011" , "011010010111111111010010100001" , "011010011000100111010010011110" , "011010011001010111010010011100" , "011010011010000111010010011001" , "011010011010101111010010010110" , "011010011011011111010010010100"
, "011010011100001111010010010001" , "011010011100111111010010001111" , "011010011101100111010010001100" , "011010011110010111010010001001" , "011010011111000111010010000111" , "011010011111110111010010000100" , "011010100000011111010010000010" , "011010100001001111010001111111" , "011010100001111111010001111100" , "011010100010100111010001111010"
, "011010100011010111010001110111" , "011010100100000111010001110101" , "011010100100110111010001110010" , "011010100101011111010001101111" , "011010100110001111010001101101" , "011010100110111111010001101010" , "011010100111100111010001100111" , "011010101000010111010001100101" , "011010101001000111010001100010" , "011010101001110111010001100000"
, "011010101010011111010001011101" , "011010101011001111010001011010" , "011010101011111111010001011000" , "011010101100100111010001010101" , "011010101101010111010001010011" , "011010101110000111010001010000" , "011010101110110111010001001101" , "011010101111011111010001001011" , "011010110000001111010001001000" , "011010110000111111010001000101"
, "011010110001100111010001000011" , "011010110010010111010001000000" , "011010110011000111010000111110" , "011010110011101111010000111011" , "011010110100011111010000111000" , "011010110101001111010000110110" , "011010110101111111010000110011" , "011010110110100111010000110000" , "011010110111010111010000101110" , "011010111000000111010000101011"
, "011010111000101111010000101000" , "011010111001011111010000100110" , "011010111010001111010000100011" , "011010111010111111010000100001" , "011010111011100111010000011110" , "011010111100010111010000011011" , "011010111101000111010000011001" , "011010111101101111010000010110" , "011010111110011111010000010011" , "011010111111001111010000010001"
, "011010111111110111010000001110" , "011011000000100111010000001011" , "011011000001010111010000001001" , "011011000001111111010000000110" , "011011000010101111010000000011" , "011011000011011111010000000001" , "011011000100001111001111111110" , "011011000100110111001111111011" , "011011000101100111001111111001" , "011011000110010111001111110110"
, "011011000110111111001111110011" , "011011000111101111001111110001" , "011011001000011111001111101110" , "011011001001000111001111101011" , "011011001001110111001111101001" , "011011001010100111001111100110" , "011011001011001111001111100011" , "011011001011111111001111100001" , "011011001100101111001111011110" , "011011001101011111001111011011"
, "011011001110000111001111011001" , "011011001110110111001111010110" , "011011001111100111001111010011" , "011011010000001111001111010001" , "011011010000111111001111001110" , "011011010001101111001111001011" , "011011010010010111001111001001" , "011011010011000111001111000110" , "011011010011110111001111000011" , "011011010100011111001111000001"
, "011011010101001111001110111110" , "011011010101111111001110111011" , "011011010110100111001110111001" , "011011010111010111001110110110" , "011011011000000111001110110011" , "011011011000101111001110110001" , "011011011001011111001110101110" , "011011011010001111001110101011" , "011011011010111111001110101000" , "011011011011100111001110100110"
, "011011011100010111001110100011" , "011011011101000111001110100000" , "011011011101101111001110011110" , "011011011110011111001110011011" , "011011011111001111001110011000" , "011011011111110111001110010110" , "011011100000100111001110010011" , "011011100001010111001110010000" , "011011100001111111001110001110" , "011011100010101111001110001011"
, "011011100011011111001110001000" , "011011100100000111001110000101" , "011011100100110111001110000011" , "011011100101100111001110000000" , "011011100110001111001101111101" , "011011100110111111001101111011" , "011011100111101111001101111000" , "011011101000010111001101110101" , "011011101001000111001101110010" , "011011101001110111001101110000"
, "011011101010011111001101101101" , "011011101011001111001101101010" , "011011101011111111001101101000" , "011011101100100111001101100101" , "011011101101010111001101100010" , "011011101110000111001101011111" , "011011101110101111001101011101" , "011011101111011111001101011010" , "011011110000001111001101010111" , "011011110000110111001101010101"
, "011011110001100111001101010010" , "011011110010010111001101001111" , "011011110010111111001101001100" , "011011110011101111001101001010" , "011011110100011111001101000111" , "011011110101000111001101000100" , "011011110101110111001101000001" , "011011110110100111001100111111" , "011011110111001111001100111100" , "011011110111111111001100111001"
, "011011111000101111001100110110" , "011011111001010111001100110100" , "011011111010000111001100110001" , "011011111010101111001100101110" , "011011111011011111001100101100" , "011011111100001111001100101001" , "011011111100110111001100100110" , "011011111101100111001100100011" , "011011111110010111001100100001" , "011011111110111111001100011110"
, "011011111111101111001100011011" , "011100000000011111001100011000" , "011100000001000111001100010110" , "011100000001110111001100010011" , "011100000010100111001100010000" , "011100000011001111001100001101" , "011100000011111111001100001011" , "011100000100101111001100001000" , "011100000101010111001100000101" , "011100000110000111001100000010"
, "011100000110110111001011111111" , "011100000111011111001011111101" , "011100001000001111001011111010" , "011100001000110111001011110111" , "011100001001100111001011110100" , "011100001010010111001011110010" , "011100001010111111001011101111" , "011100001011101111001011101100" , "011100001100011111001011101001" , "011100001101000111001011100111"
, "011100001101110111001011100100" , "011100001110100111001011100001" , "011100001111001111001011011110" , "011100001111111111001011011100" , "011100010000100111001011011001" , "011100010001010111001011010110" , "011100010010000111001011010011" , "011100010010101111001011010000" , "011100010011011111001011001110" , "011100010100001111001011001011"
, "011100010100110111001011001000" , "011100010101100111001011000101" , "011100010110010111001011000011" , "011100010110111111001011000000" , "011100010111101111001010111101" , "011100011000010111001010111010" , "011100011001000111001010110111" , "011100011001110111001010110101" , "011100011010011111001010110010" , "011100011011001111001010101111"
, "011100011011111111001010101100" , "011100011100100111001010101001" , "011100011101010111001010100111" , "011100011110000111001010100100" , "011100011110101111001010100001" , "011100011111011111001010011110" , "011100100000000111001010011011" , "011100100000110111001010011001" , "011100100001100111001010010110" , "011100100010001111001010010011"
, "011100100010111111001010010000" , "011100100011101111001010001101" , "011100100100010111001010001011" , "011100100101000111001010001000" , "011100100101101111001010000101" , "011100100110011111001010000010" , "011100100111001111001001111111" , "011100100111110111001001111101" , "011100101000100111001001111010" , "011100101001001111001001110111"
, "011100101001111111001001110100" , "011100101010101111001001110001" , "011100101011010111001001101111" , "011100101100000111001001101100" , "011100101100110111001001101001" , "011100101101011111001001100110" , "011100101110001111001001100011" , "011100101110110111001001100000" , "011100101111100111001001011110" , "011100110000010111001001011011"
, "011100110000111111001001011000" , "011100110001101111001001010101" , "011100110010010111001001010010" , "011100110011000111001001010000" , "011100110011110111001001001101" , "011100110100011111001001001010" , "011100110101001111001001000111" , "011100110101111111001001000100" , "011100110110100111001001000001" , "011100110111010111001000111111"
, "011100110111111111001000111100" , "011100111000101111001000111001" , "011100111001011111001000110110" , "011100111010000111001000110011" , "011100111010110111001000110000" , "011100111011011111001000101110" , "011100111100001111001000101011" , "011100111100111111001000101000" , "011100111101100111001000100101" , "011100111110010111001000100010"
, "011100111110111111001000011111" , "011100111111101111001000011100" , "011101000000011111001000011010" , "011101000001000111001000010111" , "011101000001110111001000010100" , "011101000010011111001000010001" , "011101000011001111001000001110" , "011101000011111111001000001011" , "011101000100100111001000001001" , "011101000101010111001000000110"
, "011101000101111111001000000011" , "011101000110101111001000000000" , "011101000111011111000111111101" , "011101001000000111000111111010" , "011101001000110111000111110111" , "011101001001011111000111110101" , "011101001010001111000111110010" , "011101001010111111000111101111" , "011101001011100111000111101100" , "011101001100010111000111101001"
, "011101001100111111000111100110" , "011101001101101111000111100011" , "011101001110011111000111100000" , "011101001111000111000111011110" , "011101001111110111000111011011" , "011101010000011111000111011000" , "011101010001001111000111010101" , "011101010001110111000111010010" , "011101010010100111000111001111" , "011101010011010111000111001100"
, "011101010011111111000111001001" , "011101010100101111000111000111" , "011101010101010111000111000100" , "011101010110000111000111000001" , "011101010110110111000110111110" , "011101010111011111000110111011" , "011101011000001111000110111000" , "011101011000110111000110110101" , "011101011001100111000110110010" , "011101011010001111000110110000"
, "011101011010111111000110101101" , "011101011011101111000110101010" , "011101011100010111000110100111" , "011101011101000111000110100100" , "011101011101101111000110100001" , "011101011110011111000110011110" , "011101011111001111000110011011" , "011101011111110111000110011000" , "011101100000100111000110010101" , "011101100001001111000110010011"
, "011101100001111111000110010000" , "011101100010100111000110001101" , "011101100011010111000110001010" , "011101100100000111000110000111" , "011101100100101111000110000100" , "011101100101011111000110000001" , "011101100110000111000101111110" , "011101100110110111000101111011" , "011101100111011111000101111000" , "011101101000001111000101110110"
, "011101101000111111000101110011" , "011101101001100111000101110000" , "011101101010010111000101101101" , "011101101010111111000101101010" , "011101101011101111000101100111" , "011101101100010111000101100100" , "011101101101000111000101100001" , "011101101101101111000101011110" , "011101101110011111000101011011" , "011101101111001111000101011000"
, "011101101111110111000101010101" , "011101110000100111000101010011" , "011101110001001111000101010000" , "011101110001111111000101001101" , "011101110010100111000101001010" , "011101110011010111000101000111" , "011101110100000111000101000100" , "011101110100101111000101000001" , "011101110101011111000100111110" , "011101110110000111000100111011"
, "011101110110110111000100111000" , "011101110111011111000100110101" , "011101111000001111000100110010" , "011101111000110111000100101111" , "011101111001100111000100101101" , "011101111010010111000100101010" , "011101111010111111000100100111" , "011101111011101111000100100100" , "011101111100010111000100100001" , "011101111101000111000100011110"
, "011101111101101111000100011011" , "011101111110011111000100011000" , "011101111111000111000100010101" , "011101111111110111000100010010" , "011110000000100111000100001111" , "011110000001001111000100001100" , "011110000001111111000100001001" , "011110000010100111000100000110" , "011110000011010111000100000011" , "011110000011111111000100000000"
, "011110000100101111000011111101" , "011110000101010111000011111010" , "011110000110000111000011111000" , "011110000110101111000011110101" , "011110000111011111000011110010" , "011110001000001111000011101111" , "011110001000110111000011101100" , "011110001001100111000011101001" , "011110001010001111000011100110" , "011110001010111111000011100011"
, "011110001011100111000011100000" , "011110001100010111000011011101" , "011110001100111111000011011010" , "011110001101101111000011010111" , "011110001110010111000011010100" , "011110001111000111000011010001" , "011110001111110111000011001110" , "011110010000011111000011001011" , "011110010001001111000011001000" , "011110010001110111000011000101"
, "011110010010100111000011000010" , "011110010011001111000010111111" , "011110010011111111000010111100" , "011110010100100111000010111001" , "011110010101010111000010110110" , "011110010101111111000010110011" , "011110010110101111000010110000" , "011110010111010111000010101101" , "011110011000000111000010101010" , "011110011000101111000010100111"
, "011110011001011111000010100100" , "011110011010000111000010100001" , "011110011010110111000010011110" , "011110011011100111000010011011" , "011110011100001111000010011000" , "011110011100111111000010010101" , "011110011101100111000010010010" , "011110011110010111000010001111" , "011110011110111111000010001100" , "011110011111101111000010001001"
, "011110100000010111000010000110" , "011110100001000111000010000011" , "011110100001101111000010000000" , "011110100010011111000001111101" , "011110100011000111000001111010" , "011110100011110111000001110111" , "011110100100011111000001110100" , "011110100101001111000001110001" , "011110100101110111000001101110" , "011110100110100111000001101011"
, "011110100111001111000001101000" , "011110100111111111000001100101" , "011110101000100111000001100010" , "011110101001010111000001011111" , "011110101010000111000001011100" , "011110101010101111000001011001" , "011110101011011111000001010110" , "011110101100000111000001010011" , "011110101100110111000001010000" , "011110101101011111000001001101"
, "011110101110001111000001001010" , "011110101110110111000001000111" , "011110101111100111000001000100" , "011110110000001111000001000001" , "011110110000111111000000111110" , "011110110001100111000000111011" , "011110110010010111000000111000" , "011110110010111111000000110101" , "011110110011101111000000110010" , "011110110100010111000000101111"
, "011110110101000111000000101100" , "011110110101101111000000101001" , "011110110110011111000000100110" , "011110110111000111000000100011" , "011110110111110111000000100000" , "011110111000011111000000011101" , "011110111001001111000000011010" , "011110111001110111000000010111" , "011110111010100111000000010100" , "011110111011001111000000010001"
, "011110111011111111000000001110" , "011110111100100111000000001011" , "011110111101010111000000001000" , "011110111101111111000000000101" , "011110111110101111000000000010" , "011110111111010110111111111111" , "011111000000000110111111111100" , "011111000000101110111111111001" , "011111000001011110111111110110" , "011111000010000110111111110010"
, "011111000010110110111111101111" , "011111000011011110111111101100" , "011111000100001110111111101001" , "011111000100110110111111100110" , "011111000101100110111111100011" , "011111000110001110111111100000" , "011111000110111110111111011101" , "011111000111100110111111011010" , "011111001000010110111111010111" , "011111001000111110111111010100"
, "011111001001101110111111010001" , "011111001010010110111111001110" , "011111001011000110111111001011" , "011111001011101110111111001000" , "011111001100011110111111000101" , "011111001101000110111111000010" , "011111001101110110111110111111" , "011111001110011110111110111011" , "011111001111000110111110111000" , "011111001111110110111110110101"
, "011111010000011110111110110010" , "011111010001001110111110101111" , "011111010001110110111110101100" , "011111010010100110111110101001" , "011111010011001110111110100110" , "011111010011111110111110100011" , "011111010100100110111110100000" , "011111010101010110111110011101" , "011111010101111110111110011010" , "011111010110101110111110010111"
, "011111010111010110111110010100" , "011111011000000110111110010000" , "011111011000101110111110001101" , "011111011001011110111110001010" , "011111011010000110111110000111" , "011111011010110110111110000100" , "011111011011011110111110000001" , "011111011100001110111101111110" , "011111011100110110111101111011" , "011111011101100110111101111000"
, "011111011110001110111101110101" , "011111011110110110111101110010" , "011111011111100110111101101110" , "011111100000001110111101101011" , "011111100000111110111101101000" , "011111100001100110111101100101" , "011111100010010110111101100010" , "011111100010111110111101011111" , "011111100011101110111101011100" , "011111100100010110111101011001"
, "011111100101000110111101010110" , "011111100101101110111101010011" , "011111100110011110111101010000" , "011111100111000110111101001100" , "011111100111110110111101001001" , "011111101000011110111101000110" , "011111101001000110111101000011" , "011111101001110110111101000000" , "011111101010011110111100111101" , "011111101011001110111100111010"
, "011111101011110110111100110111" , "011111101100100110111100110100" , "011111101101001110111100110000" , "011111101101111110111100101101" , "011111101110100110111100101010" , "011111101111010110111100100111" , "011111101111111110111100100100" , "011111110000101110111100100001" , "011111110001010110111100011110" , "011111110001111110111100011011"
, "011111110010101110111100011000" , "011111110011010110111100010100" , "011111110100000110111100010001" , "011111110100101110111100001110" , "011111110101011110111100001011" , "011111110110000110111100001000" , "011111110110110110111100000101" , "011111110111011110111100000010" , "011111111000000110111011111111" , "011111111000110110111011111011"
, "011111111001011110111011111000" , "011111111010001110111011110101" , "011111111010110110111011110010" , "011111111011100110111011101111" , "011111111100001110111011101100" , "011111111100111110111011101001" , "011111111101100110111011100101" , "011111111110001110111011100010" , "011111111110111110111011011111" , "011111111111100110111011011100"
, "100000000000010110111011011001" , "100000000000111110111011010110" , "100000000001101110111011010011" , "100000000010010110111011001111" , "100000000011000110111011001100" , "100000000011101110111011001001" , "100000000100010110111011000110" , "100000000101000110111011000011" , "100000000101101110111011000000" , "100000000110011110111010111101"
, "100000000111000110111010111001" , "100000000111110110111010110110" , "100000001000011110111010110011" , "100000001001000110111010110000" , "100000001001110110111010101101" , "100000001010011110111010101010" , "100000001011001110111010100110" , "100000001011110110111010100011" , "100000001100100110111010100000" , "100000001101001110111010011101"
, "100000001101111110111010011010" , "100000001110100110111010010111" , "100000001111001110111010010011" , "100000001111111110111010010000" , "100000010000100110111010001101" , "100000010001010110111010001010" , "100000010001111110111010000111" , "100000010010101110111010000100" , "100000010011010110111010000000" , "100000010011111110111001111101"
, "100000010100101110111001111010" , "100000010101010110111001110111" , "100000010110000110111001110100" , "100000010110101110111001110001" , "100000010111010110111001101101" , "100000011000000110111001101010" , "100000011000101110111001100111" , "100000011001011110111001100100" , "100000011010000110111001100001" , "100000011010110110111001011110"
, "100000011011011110111001011010" , "100000011100000110111001010111" , "100000011100110110111001010100" , "100000011101011110111001010001" , "100000011110001110111001001110" , "100000011110110110111001001010" , "100000011111011110111001000111" , "100000100000001110111001000100" , "100000100000110110111001000001" , "100000100001100110111000111110"
, "100000100010001110111000111010" , "100000100010111110111000110111" , "100000100011100110111000110100" , "100000100100001110111000110001" , "100000100100111110111000101110" , "100000100101100110111000101010" , "100000100110010110111000100111" , "100000100110111110111000100100" , "100000100111100110111000100001" , "100000101000010110111000011110"
, "100000101000111110111000011010" , "100000101001101110111000010111" , "100000101010010110111000010100" , "100000101010111110111000010001" , "100000101011101110111000001110" , "100000101100010110111000001010" , "100000101101000110111000000111" , "100000101101101110111000000100" , "100000101110010110111000000001" , "100000101111000110110111111110"
, "100000101111101110110111111010" , "100000110000011110110111110111" , "100000110001000110110111110100" , "100000110001101110110111110001" , "100000110010011110110111101110" , "100000110011000110110111101010" , "100000110011110110110111100111" , "100000110100011110110111100100" , "100000110101000110110111100001" , "100000110101110110110111011101"
, "100000110110011110110111011010" , "100000110111001110110111010111" , "100000110111110110110111010100" , "100000111000011110110111010001" , "100000111001001110110111001101" , "100000111001110110110111001010" , "100000111010100110110111000111" , "100000111011001110110111000100" , "100000111011110110110111000000" , "100000111100100110110110111101"
, "100000111101001110110110111010" , "100000111101110110110110110111" , "100000111110100110110110110011" , "100000111111001110110110110000" , "100000111111111110110110101101" , "100001000000100110110110101010" , "100001000001001110110110100110" , "100001000001111110110110100011" , "100001000010100110110110100000" , "100001000011010110110110011101"
, "100001000011111110110110011001" , "100001000100100110110110010110" , "100001000101010110110110010011" , "100001000101111110110110010000" , "100001000110100110110110001100" , "100001000111010110110110001001" , "100001000111111110110110000110" , "100001001000101110110110000011" , "100001001001010110110101111111" , "100001001001111110110101111100"
, "100001001010101110110101111001" , "100001001011010110110101110110" , "100001001011111110110101110010" , "100001001100101110110101101111" , "100001001101010110110101101100" , "100001001110000110110101101001" , "100001001110101110110101100101" , "100001001111010110110101100010" , "100001010000000110110101011111" , "100001010000101110110101011100"
, "100001010001010110110101011000" , "100001010010000110110101010101" , "100001010010101110110101010010" , "100001010011010110110101001111" , "100001010100000110110101001011" , "100001010100101110110101001000" , "100001010101011110110101000101" , "100001010110000110110101000001" , "100001010110101110110100111110" , "100001010111011110110100111011"
, "100001011000000110110100111000" , "100001011000101110110100110100" , "100001011001011110110100110001" , "100001011010000110110100101110" , "100001011010101110110100101011" , "100001011011011110110100100111" , "100001011100000110110100100100" , "100001011100110110110100100001" , "100001011101011110110100011101" , "100001011110000110110100011010"
, "100001011110110110110100010111" , "100001011111011110110100010100" , "100001100000000110110100010000" , "100001100000110110110100001101" , "100001100001011110110100001010" , "100001100010000110110100000110" , "100001100010110110110100000011" , "100001100011011110110100000000" , "100001100100000110110011111101" , "100001100100110110110011111001"
, "100001100101011110110011110110" , "100001100110000110110011110011" , "100001100110110110110011101111" , "100001100111011110110011101100" , "100001101000000110110011101001" , "100001101000110110110011100101" , "100001101001011110110011100010" , "100001101010001110110011011111" , "100001101010110110110011011100" , "100001101011011110110011011000"
, "100001101100001110110011010101" , "100001101100110110110011010010" , "100001101101011110110011001110" , "100001101110001110110011001011" , "100001101110110110110011001000" , "100001101111011110110011000100" , "100001110000001110110011000001" , "100001110000110110110010111110" , "100001110001011110110010111010" , "100001110010001110110010110111"
, "100001110010110110110010110100" , "100001110011011110110010110000" , "100001110100001110110010101101" , "100001110100110110110010101010" , "100001110101011110110010100110" , "100001110110001110110010100011" , "100001110110110110110010100000" , "100001110111011110110010011101" , "100001111000001110110010011001" , "100001111000110110110010010110"
, "100001111001011110110010010011" , "100001111010001110110010001111" , "100001111010110110110010001100" , "100001111011011110110010001001" , "100001111100001110110010000101" , "100001111100110110110010000010" , "100001111101011110110001111111" , "100001111110001110110001111011" , "100001111110110110110001111000" , "100001111111011110110001110101"
, "100010000000001110110001110001" , "100010000000110110110001101110" , "100010000001011110110001101011" , "100010000010001110110001100111" , "100010000010110110110001100100" , "100010000011011110110001100001" , "100010000100000110110001011101" , "100010000100110110110001011010" , "100010000101011110110001010110" , "100010000110000110110001010011"
, "100010000110110110110001010000" , "100010000111011110110001001100" , "100010001000000110110001001001" , "100010001000110110110001000110" , "100010001001011110110001000010" , "100010001010000110110000111111" , "100010001010110110110000111100" , "100010001011011110110000111000" , "100010001100000110110000110101" , "100010001100110110110000110010"
, "100010001101011110110000101110" , "100010001110000110110000101011" , "100010001110101110110000101000" , "100010001111011110110000100100" , "100010010000000110110000100001" , "100010010000101110110000011101" , "100010010001011110110000011010" , "100010010010000110110000010111" , "100010010010101110110000010011" , "100010010011011110110000010000"
, "100010010100000110110000001101" , "100010010100101110110000001001" , "100010010101011110110000000110" , "100010010110000110110000000010" , "100010010110101110101111111111" , "100010010111010110101111111100" , "100010011000000110101111111000" , "100010011000101110101111110101" , "100010011001010110101111110010" , "100010011010000110101111101110"
, "100010011010101110101111101011" , "100010011011010110101111100111" , "100010011100000110101111100100" , "100010011100101110101111100001" , "100010011101010110101111011101" , "100010011101111110101111011010" , "100010011110101110101111010111" , "100010011111010110101111010011" , "100010011111111110101111010000" , "100010100000101110101111001100"
, "100010100001010110101111001001" , "100010100001111110101111000110" , "100010100010100110101111000010" , "100010100011010110101110111111" , "100010100011111110101110111011" , "100010100100100110101110111000" , "100010100101010110101110110101" , "100010100101111110101110110001" , "100010100110100110101110101110" , "100010100111001110101110101010"
, "100010100111111110101110100111" , "100010101000100110101110100100" , "100010101001001110101110100000" , "100010101001111110101110011101" , "100010101010100110101110011001" , "100010101011001110101110010110" , "100010101011110110101110010011" , "100010101100100110101110001111" , "100010101101001110101110001100" , "100010101101110110101110001000"
, "100010101110100110101110000101" , "100010101111001110101110000010" , "100010101111110110101101111110" , "100010110000011110101101111011" , "100010110001001110101101110111" , "100010110001110110101101110100" , "100010110010011110101101110001" , "100010110011001110101101101101" , "100010110011110110101101101010" , "100010110100011110101101100110"
, "100010110101000110101101100011" , "100010110101110110101101011111" , "100010110110011110101101011100" , "100010110111000110101101011001" , "100010110111101110101101010101" , "100010111000011110101101010010" , "100010111001000110101101001110" , "100010111001101110101101001011" , "100010111010010110101101001000" , "100010111011000110101101000100"
, "100010111011101110101101000001" , "100010111100010110101100111101" , "100010111101000110101100111010" , "100010111101101110101100110110" , "100010111110010110101100110011" , "100010111110111110101100110000" , "100010111111101110101100101100" , "100011000000010110101100101001" , "100011000000111110101100100101" , "100011000001100110101100100010"
, "100011000010010110101100011110" , "100011000010111110101100011011" , "100011000011100110101100010111" , "100011000100001110101100010100" , "100011000100111110101100010001" , "100011000101100110101100001101" , "100011000110001110101100001010" , "100011000110110110101100000110" , "100011000111100110101100000011" , "100011001000001110101011111111"
, "100011001000110110101011111100" , "100011001001011110101011111000" , "100011001010001110101011110101" , "100011001010110110101011110010" , "100011001011011110101011101110" , "100011001100000110101011101011" , "100011001100110110101011100111" , "100011001101011110101011100100" , "100011001110000110101011100000" , "100011001110101110101011011101"
, "100011001111011110101011011001" , "100011010000000110101011010110" , "100011010000101110101011010010" , "100011010001010110101011001111" , "100011010010000110101011001011" , "100011010010101110101011001000" , "100011010011010110101011000101" , "100011010011111110101011000001" , "100011010100101110101010111110" , "100011010101010110101010111010"
, "100011010101111110101010110111" , "100011010110100110101010110011" , "100011010111010110101010110000" , "100011010111111110101010101100" , "100011011000100110101010101001" , "100011011001001110101010100101" , "100011011001110110101010100010" , "100011011010100110101010011110" , "100011011011001110101010011011" , "100011011011110110101010010111"
, "100011011100011110101010010100" , "100011011101001110101010010000" , "100011011101110110101010001101" , "100011011110011110101010001001" , "100011011111000110101010000110" , "100011011111110110101010000011" , "100011100000011110101001111111" , "100011100001000110101001111100" , "100011100001101110101001111000" , "100011100010010110101001110101"
, "100011100011000110101001110001" , "100011100011101110101001101110" , "100011100100010110101001101010" , "100011100100111110101001100111" , "100011100101101110101001100011" , "100011100110010110101001100000" , "100011100110111110101001011100" , "100011100111100110101001011001" , "100011101000001110101001010101" , "100011101000111110101001010010"
, "100011101001100110101001001110" , "100011101010001110101001001011" , "100011101010110110101001000111" , "100011101011100110101001000100" , "100011101100001110101001000000" , "100011101100110110101000111101" , "100011101101011110101000111001" , "100011101110000110101000110110" , "100011101110110110101000110010" , "100011101111011110101000101111"
, "100011110000000110101000101011" , "100011110000101110101000101000" , "100011110001010110101000100100" , "100011110010000110101000100001" , "100011110010101110101000011101" , "100011110011010110101000011010" , "100011110011111110101000010110" , "100011110100101110101000010010" , "100011110101010110101000001111" , "100011110101111110101000001011"
, "100011110110100110101000001000" , "100011110111001110101000000100" , "100011110111111110101000000001" , "100011111000100110100111111101" , "100011111001001110100111111010" , "100011111001110110100111110110" , "100011111010011110100111110011" , "100011111011001110100111101111" , "100011111011110110100111101100" , "100011111100011110100111101000"
, "100011111101000110100111100101" , "100011111101101110100111100001" , "100011111110011110100111011110" , "100011111111000110100111011010" , "100011111111101110100111010111" , "100100000000010110100111010011" , "100100000000111110100111010000" , "100100000001101110100111001100" , "100100000010010110100111001000" , "100100000010111110100111000101"
, "100100000011100110100111000001" , "100100000100001110100110111110" , "100100000100110110100110111010" , "100100000101100110100110110111" , "100100000110001110100110110011" , "100100000110110110100110110000" , "100100000111011110100110101100" , "100100001000000110100110101001" , "100100001000110110100110100101" , "100100001001011110100110100001"
, "100100001010000110100110011110" , "100100001010101110100110011010" , "100100001011010110100110010111" , "100100001100000110100110010011" , "100100001100101110100110010000" , "100100001101010110100110001100" , "100100001101111110100110001001" , "100100001110100110100110000101" , "100100001111001110100110000001" , "100100001111111110100101111110"
, "100100010000100110100101111010" , "100100010001001110100101110111" , "100100010001110110100101110011" , "100100010010011110100101110000" , "100100010011001110100101101100" , "100100010011110110100101101001" , "100100010100011110100101100101" , "100100010101000110100101100001" , "100100010101101110100101011110" , "100100010110010110100101011010"
, "100100010111000110100101010111" , "100100010111101110100101010011" , "100100011000010110100101010000" , "100100011000111110100101001100" , "100100011001100110100101001000" , "100100011010001110100101000101" , "100100011010111110100101000001" , "100100011011100110100100111110" , "100100011100001110100100111010" , "100100011100110110100100110111"
, "100100011101011110100100110011" , "100100011110000110100100101111" , "100100011110110110100100101100" , "100100011111011110100100101000" , "100100100000000110100100100101" , "100100100000101110100100100001" , "100100100001010110100100011101" , "100100100001111110100100011010" , "100100100010101110100100010110" , "100100100011010110100100010011"
, "100100100011111110100100001111" , "100100100100100110100100001100" , "100100100101001110100100001000" , "100100100101110110100100000100" , "100100100110011110100100000001" , "100100100111001110100011111101" , "100100100111110110100011111010" , "100100101000011110100011110110" , "100100101001000110100011110010" , "100100101001101110100011101111"
, "100100101010010110100011101011" , "100100101011000110100011101000" , "100100101011101110100011100100" , "100100101100010110100011100000" , "100100101100111110100011011101" , "100100101101100110100011011001" , "100100101110001110100011010110" , "100100101110110110100011010010" , "100100101111100110100011001110" , "100100110000001110100011001011"
, "100100110000110110100011000111" , "100100110001011110100011000100" , "100100110010000110100011000000" , "100100110010101110100010111100" , "100100110011010110100010111001" , "100100110100000110100010110101" , "100100110100101110100010110001" , "100100110101010110100010101110" , "100100110101111110100010101010" , "100100110110100110100010100111"
, "100100110111001110100010100011" , "100100110111110110100010011111" , "100100111000011110100010011100" , "100100111001001110100010011000" , "100100111001110110100010010101" , "100100111010011110100010010001" , "100100111011000110100010001101" , "100100111011101110100010001010" , "100100111100010110100010000110" , "100100111100111110100010000010"
, "100100111101101110100001111111" , "100100111110010110100001111011" , "100100111110111110100001111000" , "100100111111100110100001110100" , "100101000000001110100001110000" , "100101000000110110100001101101" , "100101000001011110100001101001" , "100101000010000110100001100101" , "100101000010110110100001100010" , "100101000011011110100001011110"
, "100101000100000110100001011010" , "100101000100101110100001010111" , "100101000101010110100001010011" , "100101000101111110100001010000" , "100101000110100110100001001100" , "100101000111001110100001001000" , "100101000111111110100001000101" , "100101001000100110100001000001" , "100101001001001110100000111101" , "100101001001110110100000111010"
, "100101001010011110100000110110" , "100101001011000110100000110010" , "100101001011101110100000101111" , "100101001100010110100000101011" , "100101001100111110100000100111" , "100101001101101110100000100100" , "100101001110010110100000100000" , "100101001110111110100000011100" , "100101001111100110100000011001" , "100101010000001110100000010101"
, "100101010000110110100000010001" , "100101010001011110100000001110" , "100101010010000110100000001010" , "100101010010101110100000000110" , "100101010011011110100000000011" , "100101010100000110011111111111" , "100101010100101110011111111011" , "100101010101010110011111111000" , "100101010101111110011111110100" , "100101010110100110011111110000"
, "100101010111001110011111101101" , "100101010111110110011111101001" , "100101011000011110011111100101" , "100101011001000110011111100010" , "100101011001110110011111011110" , "100101011010011110011111011010" , "100101011011000110011111010111" , "100101011011101110011111010011" , "100101011100010110011111001111" , "100101011100111110011111001100"
, "100101011101100110011111001000" , "100101011110001110011111000100" , "100101011110110110011111000001" , "100101011111011110011110111101" , "100101100000001110011110111001" , "100101100000110110011110110110" , "100101100001011110011110110010" , "100101100010000110011110101110" , "100101100010101110011110101011" , "100101100011010110011110100111"
, "100101100011111110011110100011" , "100101100100100110011110100000" , "100101100101001110011110011100" , "100101100101110110011110011000" , "100101100110011110011110010101" , "100101100111000110011110010001" , "100101100111110110011110001101" , "100101101000011110011110001001" , "100101101001000110011110000110" , "100101101001101110011110000010"
, "100101101010010110011101111110" , "100101101010111110011101111011" , "100101101011100110011101110111" , "100101101100001110011101110011" , "100101101100110110011101110000" , "100101101101011110011101101100" , "100101101110000110011101101000" , "100101101110101110011101100100" , "100101101111011110011101100001" , "100101110000000110011101011101"
, "100101110000101110011101011001" , "100101110001010110011101010110" , "100101110001111110011101010010" , "100101110010100110011101001110" , "100101110011001110011101001010" , "100101110011110110011101000111" , "100101110100011110011101000011" , "100101110101000110011100111111" , "100101110101101110011100111100" , "100101110110010110011100111000"
, "100101110110111110011100110100" , "100101110111100110011100110000" , "100101111000001110011100101101" , "100101111000111110011100101001" , "100101111001100110011100100101" , "100101111010001110011100100010" , "100101111010110110011100011110" , "100101111011011110011100011010" , "100101111100000110011100010110" , "100101111100101110011100010011"
, "100101111101010110011100001111" , "100101111101111110011100001011" , "100101111110100110011100001000" , "100101111111001110011100000100" , "100101111111110110011100000000" , "100110000000011110011011111100" , "100110000001000110011011111001" , "100110000001101110011011110101" , "100110000010010110011011110001" , "100110000010111110011011101101"
, "100110000011101110011011101010" , "100110000100010110011011100110" , "100110000100111110011011100010" , "100110000101100110011011011110" , "100110000110001110011011011011" , "100110000110110110011011010111" , "100110000111011110011011010011" , "100110001000000110011011010000" , "100110001000101110011011001100" , "100110001001010110011011001000"
, "100110001001111110011011000100" , "100110001010100110011011000001" , "100110001011001110011010111101" , "100110001011110110011010111001" , "100110001100011110011010110101" , "100110001101000110011010110010" , "100110001101101110011010101110" , "100110001110010110011010101010" , "100110001110111110011010100110" , "100110001111100110011010100011"
, "100110010000001110011010011111" , "100110010000110110011010011011" , "100110010001011110011010010111" , "100110010010001110011010010011" , "100110010010110110011010010000" , "100110010011011110011010001100" , "100110010100000110011010001000" , "100110010100101110011010000100" , "100110010101010110011010000001" , "100110010101111110011001111101"
, "100110010110100110011001111001" , "100110010111001110011001110101" , "100110010111110110011001110010" , "100110011000011110011001101110" , "100110011001000110011001101010" , "100110011001101110011001100110" , "100110011010010110011001100011" , "100110011010111110011001011111" , "100110011011100110011001011011" , "100110011100001110011001010111"
, "100110011100110110011001010011" , "100110011101011110011001010000" , "100110011110000110011001001100" , "100110011110101110011001001000" , "100110011111010110011001000100" , "100110011111111110011001000001" , "100110100000100110011000111101" , "100110100001001110011000111001" , "100110100001110110011000110101" , "100110100010011110011000110001"
, "100110100011000110011000101110" , "100110100011101110011000101010" , "100110100100010110011000100110" , "100110100100111110011000100010" , "100110100101100110011000011111" , "100110100110001110011000011011" , "100110100110110110011000010111" , "100110100111011110011000010011" , "100110101000000110011000001111" , "100110101000101110011000001100"
, "100110101001010110011000001000" , "100110101001111110011000000100" , "100110101010100110011000000000" , "100110101011001110010111111100" , "100110101011110110010111111001" , "100110101100011110010111110101" , "100110101101000110010111110001" , "100110101101101110010111101101" , "100110101110010110010111101001" , "100110101110111110010111100110"
, "100110101111100110010111100010" , "100110110000001110010111011110" , "100110110000110110010111011010" , "100110110001011110010111010110" , "100110110010000110010111010011" , "100110110010101110010111001111" , "100110110011010110010111001011" , "100110110011111110010111000111" , "100110110100100110010111000011" , "100110110101001110010111000000"
, "100110110101110110010110111100" , "100110110110011110010110111000" , "100110110111000110010110110100" , "100110110111101110010110110000" , "100110111000010110010110101100" , "100110111000111110010110101001" , "100110111001100110010110100101" , "100110111010001110010110100001" , "100110111010110110010110011101" , "100110111011011110010110011001"
, "100110111100000110010110010110" , "100110111100101110010110010010" , "100110111101010110010110001110" , "100110111101111110010110001010" , "100110111110100110010110000110" , "100110111111001110010110000010" , "100110111111110110010101111111" , "100111000000011110010101111011" , "100111000001000110010101110111" , "100111000001101110010101110011"
, "100111000010010110010101101111" , "100111000010111110010101101011" , "100111000011100110010101101000" , "100111000100001110010101100100" , "100111000100110110010101100000" , "100111000101011110010101011100" , "100111000110000110010101011000" , "100111000110101110010101010100" , "100111000111010110010101010001" , "100111000111111110010101001101"
, "100111001000100110010101001001" , "100111001001001110010101000101" , "100111001001110110010101000001" , "100111001010011110010100111101" , "100111001011000110010100111010" , "100111001011101110010100110110" , "100111001100010110010100110010" , "100111001100111110010100101110" , "100111001101100110010100101010" , "100111001110001110010100100110"
, "100111001110110110010100100010" , "100111001111010110010100011111" , "100111001111111110010100011011" , "100111010000100110010100010111" , "100111010001001110010100010011" , "100111010001110110010100001111" , "100111010010011110010100001011" , "100111010011000110010100000111" , "100111010011101110010100000100" , "100111010100010110010100000000"
, "100111010100111110010011111100" , "100111010101100110010011111000" , "100111010110001110010011110100" , "100111010110110110010011110000" , "100111010111011110010011101100" , "100111011000000110010011101001" , "100111011000101110010011100101" , "100111011001010110010011100001" , "100111011001111110010011011101" , "100111011010100110010011011001"
, "100111011011001110010011010101" , "100111011011110110010011010001" , "100111011100011110010011001101" , "100111011101000110010011001010" , "100111011101100110010011000110" , "100111011110001110010011000010" , "100111011110110110010010111110" , "100111011111011110010010111010" , "100111100000000110010010110110" , "100111100000101110010010110010"
, "100111100001010110010010101110" , "100111100001111110010010101011" , "100111100010100110010010100111" , "100111100011001110010010100011" , "100111100011110110010010011111" , "100111100100011110010010011011" , "100111100101000110010010010111" , "100111100101101110010010010011" , "100111100110010110010010001111" , "100111100110111110010010001011"
, "100111100111100110010010001000" , "100111101000000110010010000100" , "100111101000101110010010000000" , "100111101001010110010001111100" , "100111101001111110010001111000" , "100111101010100110010001110100" , "100111101011001110010001110000" , "100111101011110110010001101100" , "100111101100011110010001101000" , "100111101101000110010001100101"
, "100111101101101110010001100001" , "100111101110010110010001011101" , "100111101110111110010001011001" , "100111101111100110010001010101" , "100111110000001110010001010001" , "100111110000101110010001001101" , "100111110001010110010001001001" , "100111110001111110010001000101" , "100111110010100110010001000001" , "100111110011001110010000111110"
, "100111110011110110010000111010" , "100111110100011110010000110110" , "100111110101000110010000110010" , "100111110101101110010000101110" , "100111110110010110010000101010" , "100111110110111110010000100110" , "100111110111100110010000100010" , "100111111000000110010000011110" , "100111111000101110010000011010" , "100111111001010110010000010110"
, "100111111001111110010000010010" , "100111111010100110010000001111" , "100111111011001110010000001011" , "100111111011110110010000000111" , "100111111100011110010000000011" , "100111111101000110001111111111" , "100111111101101110001111111011" , "100111111110010110001111110111" , "100111111110110110001111110011" , "100111111111011110001111101111"
, "101000000000000110001111101011" , "101000000000101110001111100111" , "101000000001010110001111100011" , "101000000001111110001111011111" , "101000000010100110001111011100" , "101000000011001110001111011000" , "101000000011110110001111010100" , "101000000100011110001111010000" , "101000000101000110001111001100" , "101000000101100110001111001000"
, "101000000110001110001111000100" , "101000000110110110001111000000" , "101000000111011110001110111100" , "101000001000000110001110111000" , "101000001000101110001110110100" , "101000001001010110001110110000" , "101000001001111110001110101100" , "101000001010100110001110101000" , "101000001011000110001110100100" , "101000001011101110001110100000"
, "101000001100010110001110011101" , "101000001100111110001110011001" , "101000001101100110001110010101" , "101000001110001110001110010001" , "101000001110110110001110001101" , "101000001111011110001110001001" , "101000010000000110001110000101" , "101000010000100110001110000001" , "101000010001001110001101111101" , "101000010001110110001101111001"
, "101000010010011110001101110101" , "101000010011000110001101110001" , "101000010011101110001101101101" , "101000010100010110001101101001" , "101000010100111110001101100101" , "101000010101100110001101100001" , "101000010110000110001101011101" , "101000010110101110001101011001" , "101000010111010110001101010101" , "101000010111111110001101010001"
, "101000011000100110001101001101" , "101000011001001110001101001001" , "101000011001110110001101000110" , "101000011010011110001101000010" , "101000011010111110001100111110" , "101000011011100110001100111010" , "101000011100001110001100110110" , "101000011100110110001100110010" , "101000011101011110001100101110" , "101000011110000110001100101010"
, "101000011110101110001100100110" , "101000011111001110001100100010" , "101000011111110110001100011110" , "101000100000011110001100011010" , "101000100001000110001100010110" , "101000100001101110001100010010" , "101000100010010110001100001110" , "101000100010111110001100001010" , "101000100011100110001100000110" , "101000100100000110001100000010"
, "101000100100101110001011111110" , "101000100101010110001011111010" , "101000100101111110001011110110" , "101000100110100110001011110010" , "101000100111001110001011101110" , "101000100111110110001011101010" , "101000101000010110001011100110" , "101000101000111110001011100010" , "101000101001100110001011011110" , "101000101010001110001011011010"
, "101000101010110110001011010110" , "101000101011011110001011010010" , "101000101011111110001011001110" , "101000101100100110001011001010" , "101000101101001110001011000110" , "101000101101110110001011000010" , "101000101110011110001010111110" , "101000101111000110001010111010" , "101000101111101110001010110110" , "101000110000001110001010110010"
, "101000110000110110001010101110" , "101000110001011110001010101010" , "101000110010000110001010100110" , "101000110010101110001010100010" , "101000110011010110001010011110" , "101000110011110110001010011010" , "101000110100011110001010010110" , "101000110101000110001010010010" , "101000110101101110001010001110" , "101000110110010110001010001010"
, "101000110110111110001010000110" , "101000110111011110001010000010" , "101000111000000110001001111110" , "101000111000101110001001111010" , "101000111001010110001001110110" , "101000111001111110001001110010" , "101000111010100110001001101110" , "101000111011000110001001101010" , "101000111011101110001001100110" , "101000111100010110001001100010"
, "101000111100111110001001011110" , "101000111101100110001001011010" , "101000111110001110001001010110" , "101000111110101110001001010010" , "101000111111010110001001001110" , "101000111111111110001001001010" , "101001000000100110001001000110" , "101001000001001110001001000010" , "101001000001110110001000111110" , "101001000010010110001000111010"
, "101001000010111110001000110110" , "101001000011100110001000110010" , "101001000100001110001000101110" , "101001000100110110001000101010" , "101001000101011110001000100110" , "101001000101111110001000100001" , "101001000110100110001000011101" , "101001000111001110001000011001" , "101001000111110110001000010101" , "101001001000011110001000010001"
, "101001001000111110001000001101" , "101001001001100110001000001001" , "101001001010001110001000000101" , "101001001010110110001000000001" , "101001001011011110000111111101" , "101001001011111110000111111001" , "101001001100100110000111110101" , "101001001101001110000111110001" , "101001001101110110000111101101" , "101001001110011110000111101001"
, "101001001110111110000111100101" , "101001001111100110000111100001" , "101001010000001110000111011101" , "101001010000110110000111011001" , "101001010001011110000111010101" , "101001010010000110000111010001" , "101001010010100110000111001101" , "101001010011001110000111001001" , "101001010011110110000111000100" , "101001010100011110000111000000"
, "101001010101000110000110111100" , "101001010101100110000110111000" , "101001010110001110000110110100" , "101001010110110110000110110000" , "101001010111011110000110101100" , "101001010111111110000110101000" , "101001011000100110000110100100" , "101001011001001110000110100000" , "101001011001110110000110011100" , "101001011010011110000110011000"
, "101001011010111110000110010100" , "101001011011100110000110010000" , "101001011100001110000110001100" , "101001011100110110000110001000" , "101001011101011110000110000011" , "101001011101111110000101111111" , "101001011110100110000101111011" , "101001011111001110000101110111" , "101001011111110110000101110011" , "101001100000011110000101101111"
, "101001100000111110000101101011" , "101001100001100110000101100111" , "101001100010001110000101100011" , "101001100010110110000101011111" , "101001100011010110000101011011" , "101001100011111110000101010111" , "101001100100100110000101010011" , "101001100101001110000101001110" , "101001100101110110000101001010" , "101001100110010110000101000110"
, "101001100110111110000101000010" , "101001100111100110000100111110" , "101001101000001110000100111010" , "101001101000101110000100110110" , "101001101001010110000100110010" , "101001101001111110000100101110" , "101001101010100110000100101010" , "101001101011000110000100100110" , "101001101011101110000100100001" , "101001101100010110000100011101"
, "101001101100111110000100011001" , "101001101101100110000100010101" , "101001101110000110000100010001" , "101001101110101110000100001101" , "101001101111010110000100001001" , "101001101111111110000100000101" , "101001110000011110000100000001" , "101001110001000110000011111101" , "101001110001101110000011111001" , "101001110010010110000011110100"
, "101001110010110110000011110000" , "101001110011011110000011101100" , "101001110100000110000011101000" , "101001110100101110000011100100" , "101001110101001110000011100000" , "101001110101110110000011011100" , "101001110110011110000011011000" , "101001110111000110000011010100" , "101001110111100110000011001111" , "101001111000001110000011001011"
, "101001111000110110000011000111" , "101001111001011110000011000011" , "101001111001111110000010111111" , "101001111010100110000010111011" , "101001111011001110000010110111" , "101001111011110110000010110011" , "101001111100010110000010101111" , "101001111100111110000010101010" , "101001111101100110000010100110" , "101001111110001110000010100010"
, "101001111110101110000010011110" , "101001111111010110000010011010" , "101001111111111110000010010110" , "101010000000100110000010010010" , "101010000001000110000010001110" , "101010000001101110000010001001" , "101010000010010110000010000101" , "101010000010111110000010000001" , "101010000011011110000001111101" , "101010000100000110000001111001"
, "101010000100101110000001110101" , "101010000101010110000001110001" , "101010000101110110000001101101" , "101010000110011110000001101000" , "101010000111000110000001100100" , "101010000111100110000001100000" , "101010001000001110000001011100" , "101010001000110110000001011000" , "101010001001011110000001010100" , "101010001001111110000001010000"
, "101010001010100110000001001011" , "101010001011001110000001000111" , "101010001011110110000001000011" , "101010001100010110000000111111" , "101010001100111110000000111011" , "101010001101100110000000110111" , "101010001110000110000000110011" , "101010001110101110000000101110" , "101010001111010110000000101010" , "101010001111111110000000100110"
, "101010010000011110000000100010" , "101010010001000110000000011110" , "101010010001101110000000011010" , "101010010010001110000000010110" , "101010010010110110000000010001" , "101010010011011110000000001101" , "101010010100000110000000001001" , "101010010100100110000000000101" , "101010010101001110000000000001" , "101010010101110101111111111101"
, "101010010110010101111111111001" , "101010010110111101111111110100" , "101010010111100101111111110000" , "101010011000001101111111101100" , "101010011000101101111111101000" , "101010011001010101111111100100" , "101010011001111101111111100000" , "101010011010011101111111011011" , "101010011011000101111111010111" , "101010011011101101111111010011"
, "101010011100010101111111001111" , "101010011100110101111111001011" , "101010011101011101111111000111" , "101010011110000101111111000010" , "101010011110100101111110111110" , "101010011111001101111110111010" , "101010011111110101111110110110" , "101010100000010101111110110010" , "101010100000111101111110101110" , "101010100001100101111110101001"
, "101010100010001101111110100101" , "101010100010101101111110100001" , "101010100011010101111110011101" , "101010100011111101111110011001" , "101010100100011101111110010100" , "101010100101000101111110010000" , "101010100101101101111110001100" , "101010100110001101111110001000" , "101010100110110101111110000100" , "101010100111011101111110000000"
, "101010100111111101111101111011" , "101010101000100101111101110111" , "101010101001001101111101110011" , "101010101001110101111101101111" , "101010101010010101111101101011" , "101010101010111101111101100110" , "101010101011100101111101100010" , "101010101100000101111101011110" , "101010101100101101111101011010" , "101010101101010101111101010110"
, "101010101101110101111101010001" , "101010101110011101111101001101" , "101010101111000101111101001001" , "101010101111100101111101000101" , "101010110000001101111101000001" , "101010110000110101111100111100" , "101010110001010101111100111000" , "101010110001111101111100110100" , "101010110010100101111100110000" , "101010110011000101111100101100"
, "101010110011101101111100100111" , "101010110100010101111100100011" , "101010110100110101111100011111" , "101010110101011101111100011011" , "101010110110000101111100010111" , "101010110110100101111100010010" , "101010110111001101111100001110" , "101010110111110101111100001010" , "101010111000010101111100000110" , "101010111000111101111100000010"
, "101010111001100101111011111101" , "101010111010000101111011111001" , "101010111010101101111011110101" , "101010111011010101111011110001" , "101010111011110101111011101101" , "101010111100011101111011101000" , "101010111101000101111011100100" , "101010111101100101111011100000" , "101010111110001101111011011100" , "101010111110110101111011010111"
, "101010111111010101111011010011" , "101010111111111101111011001111" , "101011000000100101111011001011" , "101011000001000101111011000111" , "101011000001101101111011000010" , "101011000010010101111010111110" , "101011000010110101111010111010" , "101011000011011101111010110110" , "101011000100000101111010110001" , "101011000100100101111010101101"
, "101011000101001101111010101001" , "101011000101101101111010100101" , "101011000110010101111010100001" , "101011000110111101111010011100" , "101011000111011101111010011000" , "101011001000000101111010010100" , "101011001000101101111010010000" , "101011001001001101111010001011" , "101011001001110101111010000111" , "101011001010011101111010000011"
, "101011001010111101111001111111" , "101011001011100101111001111010" , "101011001100001101111001110110" , "101011001100101101111001110010" , "101011001101010101111001101110" , "101011001101110101111001101001" , "101011001110011101111001100101" , "101011001111000101111001100001" , "101011001111100101111001011101" , "101011010000001101111001011000"
, "101011010000110101111001010100" , "101011010001010101111001010000" , "101011010001111101111001001100" , "101011010010011101111001001000" , "101011010011000101111001000011" , "101011010011101101111000111111" , "101011010100001101111000111011" , "101011010100110101111000110111" , "101011010101011101111000110010" , "101011010101111101111000101110"
, "101011010110100101111000101010" , "101011010111000101111000100101" , "101011010111101101111000100001" , "101011011000010101111000011101" , "101011011000110101111000011001" , "101011011001011101111000010100" , "101011011010000101111000010000" , "101011011010100101111000001100" , "101011011011001101111000001000" , "101011011011101101111000000011"
, "101011011100010101110111111111" , "101011011100111101110111111011" , "101011011101011101110111110111" , "101011011110000101110111110010" , "101011011110100101110111101110" , "101011011111001101110111101010" , "101011011111110101110111100110" , "101011100000010101110111100001" , "101011100000111101110111011101" , "101011100001100101110111011001"
, "101011100010000101110111010100" , "101011100010101101110111010000" , "101011100011001101110111001100" , "101011100011110101110111001000" , "101011100100011101110111000011" , "101011100100111101110110111111" , "101011100101100101110110111011" , "101011100110000101110110110111" , "101011100110101101110110110010" , "101011100111010101110110101110"
, "101011100111110101110110101010" , "101011101000011101110110100101" , "101011101000111101110110100001" , "101011101001100101110110011101" , "101011101010001101110110011001" , "101011101010101101110110010100" , "101011101011010101110110010000" , "101011101011110101110110001100" , "101011101100011101110110000111" , "101011101100111101110110000011"
, "101011101101100101110101111111" , "101011101110001101110101111010" , "101011101110101101110101110110" , "101011101111010101110101110010" , "101011101111110101110101101110" , "101011110000011101110101101001" , "101011110001000101110101100101" , "101011110001100101110101100001" , "101011110010001101110101011100" , "101011110010101101110101011000"
, "101011110011010101110101010100" , "101011110011111101110101010000" , "101011110100011101110101001011" , "101011110101000101110101000111" , "101011110101100101110101000011" , "101011110110001101110100111110" , "101011110110101101110100111010" , "101011110111010101110100110110" , "101011110111111101110100110001" , "101011111000011101110100101101"
, "101011111001000101110100101001" , "101011111001100101110100100100" , "101011111010001101110100100000" , "101011111010101101110100011100" , "101011111011010101110100011000" , "101011111011111101110100010011" , "101011111100011101110100001111" , "101011111101000101110100001011" , "101011111101100101110100000110" , "101011111110001101110100000010"
, "101011111110101101110011111110" , "101011111111010101110011111001" , "101011111111111101110011110101" , "101100000000011101110011110001" , "101100000001000101110011101100" , "101100000001100101110011101000" , "101100000010001101110011100100" , "101100000010101101110011011111" , "101100000011010101110011011011" , "101100000011110101110011010111"
, "101100000100011101110011010010" , "101100000101000101110011001110" , "101100000101100101110011001010" , "101100000110001101110011000101" , "101100000110101101110011000001" , "101100000111010101110010111101" , "101100000111110101110010111000" , "101100001000011101110010110100" , "101100001000111101110010110000" , "101100001001100101110010101011"
, "101100001010001101110010100111" , "101100001010101101110010100011" , "101100001011010101110010011110" , "101100001011110101110010011010" , "101100001100011101110010010110" , "101100001100111101110010010001" , "101100001101100101110010001101" , "101100001110000101110010001001" , "101100001110101101110010000100" , "101100001111001101110010000000"
, "101100001111110101110001111100" , "101100010000010101110001110111" , "101100010000111101110001110011" , "101100010001100101110001101111" , "101100010010000101110001101010" , "101100010010101101110001100110" , "101100010011001101110001100010" , "101100010011110101110001011101" , "101100010100010101110001011001" , "101100010100111101110001010101"
, "101100010101011101110001010000" , "101100010110000101110001001100" , "101100010110100101110001001000" , "101100010111001101110001000011" , "101100010111101101110000111111" , "101100011000010101110000111010" , "101100011000110101110000110110" , "101100011001011101110000110010" , "101100011010000101110000101101" , "101100011010100101110000101001"
, "101100011011001101110000100101" , "101100011011101101110000100000" , "101100011100010101110000011100" , "101100011100110101110000011000" , "101100011101011101110000010011" , "101100011101111101110000001111" , "101100011110100101110000001010" , "101100011111000101110000000110" , "101100011111101101110000000010" , "101100100000001101101111111101"
, "101100100000110101101111111001" , "101100100001010101101111110101" , "101100100001111101101111110000" , "101100100010011101101111101100" , "101100100011000101101111101000" , "101100100011100101101111100011" , "101100100100001101101111011111" , "101100100100101101101111011010" , "101100100101010101101111010110" , "101100100101110101101111010010"
, "101100100110011101101111001101" , "101100100110111101101111001001" , "101100100111100101101111000101" , "101100101000000101101111000000" , "101100101000101101101110111100" , "101100101001001101101110110111" , "101100101001110101101110110011" , "101100101010010101101110101111" , "101100101010111101101110101010" , "101100101011011101101110100110"
, "101100101100000101101110100001" , "101100101100100101101110011101" , "101100101101001101101110011001" , "101100101101101101101110010100" , "101100101110010101101110010000" , "101100101110110101101110001100" , "101100101111011101101110000111" , "101100101111111101101110000011" , "101100110000100101101101111110" , "101100110001000101101101111010"
, "101100110001101101101101110110" , "101100110010001101101101110001" , "101100110010110101101101101101" , "101100110011010101101101101000" , "101100110011111101101101100100" , "101100110100011101101101100000" , "101100110101000101101101011011" , "101100110101100101101101010111" , "101100110110001101101101010010" , "101100110110101101101101001110"
, "101100110111010101101101001010" , "101100110111110101101101000101" , "101100111000011101101101000001" , "101100111000111101101100111100" , "101100111001100101101100111000" , "101100111010000101101100110100" , "101100111010101101101100101111" , "101100111011001101101100101011" , "101100111011110101101100100110" , "101100111100010101101100100010"
, "101100111100110101101100011101" , "101100111101011101101100011001" , "101100111101111101101100010101" , "101100111110100101101100010000" , "101100111111000101101100001100" , "101100111111101101101100000111" , "101101000000001101101100000011" , "101101000000110101101011111111" , "101101000001010101101011111010" , "101101000001111101101011110110"
, "101101000010011101101011110001" , "101101000011000101101011101101" , "101101000011100101101011101000" , "101101000100001101101011100100" , "101101000100101101101011100000" , "101101000101001101101011011011" , "101101000101110101101011010111" , "101101000110010101101011010010" , "101101000110111101101011001110" , "101101000111011101101011001001"
, "101101001000000101101011000101" , "101101001000100101101011000001" , "101101001001001101101010111100" , "101101001001101101101010111000" , "101101001010010101101010110011" , "101101001010110101101010101111" , "101101001011010101101010101010" , "101101001011111101101010100110" , "101101001100011101101010100010" , "101101001101000101101010011101"
, "101101001101100101101010011001" , "101101001110001101101010010100" , "101101001110101101101010010000" , "101101001111010101101010001011" , "101101001111110101101010000111" , "101101010000010101101010000010"
);
end a;

