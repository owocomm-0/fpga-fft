
library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
-- read delay is 2 cycles

entity twiddleRom1024 is
	port(clk: in std_logic;
			romAddr: in unsigned(7-1 downto 0);
			romData: out std_logic_vector(30-1 downto 0)
			);
end entity;
architecture a of twiddleRom1024 is
	constant romDepthOrder: integer := 7;
	constant romDepth: integer := 2**romDepthOrder;
	constant romWidth: integer := 30;
	--ram
	type ram1t is array(0 to romDepth-1) of
		std_logic_vector(romWidth-1 downto 0);
	signal rom: ram1t;
	signal addr1: unsigned(romDepthOrder-1 downto 0) := (others=>'0');
	signal data0,data1: std_logic_vector(romWidth-1 downto 0) := (others=>'0');
begin
	addr1 <= romAddr when rising_edge(clk);
	data0 <= rom(to_integer(addr1));
	data1 <= data0 when rising_edge(clk);
	romData <= data1;
	rom <= (
"000000011001001111111111111111" , "000000110010010111111111111110" , "000001001011011111111111111010" , "000001100100100111111111110110" , "000001111101101111111111110001" , "000010010110110111111111101010" , "000010101111111111111111100010" , "000011001001000111111111011001" , "000011100010001111111111001110" , "000011111011001111111111000010"
, "000100010100010111111110110101" , "000100101101011111111110100111" , "000101000110011111111110011000" , "000101011111011111111110000111" , "000101111000100111111101110101" , "000110010001100111111101100010" , "000110101010100111111101001110" , "000111000011100111111100111000" , "000111011100100111111100100010" , "000111110101011111111100001010"
, "001000001110011111111011110000" , "001000100111010111111011010110" , "001001000000001111111010111010" , "001001011001000111111010011101" , "001001110001111111111001111111" , "001010001010101111111001100000" , "001010100011100111111000111111" , "001010111100010111111000011110" , "001011010101000111110111111011" , "001011101101110111110111010110"
, "001100000110011111110110110001" , "001100011111001111110110001010" , "001100110111110111110101100011" , "001101010000011111110100111010" , "001101101000111111110100001111" , "001110000001100111110011100100" , "001110011010000111110010110111" , "001110110010011111110010001001" , "001111001010111111110001011010" , "001111100011010111110000101010"
, "001111111011101111101111111001" , "010000010011111111101111000110" , "010000101100010111101110010010" , "010001000100100111101101011101" , "010001011100101111101100100111" , "010001110100111111101011101111" , "010010001100111111101010110111" , "010010100101000111101001111101" , "010010111101000111101001000010" , "010011010101000111101000000110"
, "010011101101000111100111001001" , "010100000100111111100110001010" , "010100011100101111100101001010" , "010100110100100111100100001010" , "010101001100010111100011001000" , "010101100011111111100010000101" , "010101111011100111100001000000" , "010110010011001111011111111011" , "010110101010101111011110110100" , "010111000010001111011101101100"
, "010111011001100111011100100011" , "010111110000111111011011011001" , "011000001000010111011010001110" , "011000011111100111011001000010" , "011000110110101111010111110100" , "011001001101110111010110100110" , "011001100100111111010101010110" , "011001111011111111010100000101" , "011010010010111111010010110011" , "011010101001110111010001100000"
, "011011000000100111010000001011" , "011011010111010111001110110110" , "011011101110000111001101011111" , "011100000100101111001100001000" , "011100011011001111001010101111" , "011100110001101111001001010101" , "011101001000000111000111111010" , "011101011110011111000110011110" , "011101110100101111000101000001" , "011110001010111111000011100011"
, "011110100001000111000010000011" , "011110110111000111000000100011" , "011111001101000110111111000010" , "011111100010111110111101011111" , "011111111000110110111011111011" , "100000001110100110111010010111" , "100000100100001110111000110001" , "100000111001110110110111001010" , "100001001111010110110101100010" , "100001100100110110110011111001"
, "100001111010001110110010001111" , "100010001111011110110000100100" , "100010100100100110101110111000" , "100010111001101110101101001011" , "100011001110101110101011011101" , "100011100011101110101001101110" , "100011111000100110100111111101" , "100100001101010110100110001100" , "100100100001111110100100011010" , "100100110110100110100010100111"
, "100101001011000110100000110010" , "100101011111011110011110111101" , "100101110011110110011101000111" , "100110001000000110011011010000" , "100110011100001110011001010111" , "100110110000001110010111011110" , "100111000100001110010101100100" , "100111011000000110010011101001" , "100111101011110110010001101100" , "100111111111011110001111101111"
, "101000010011000110001101110001" , "101000100110100110001011110010" , "101000111001111110001001110010" , "101001001101001110000111110001" , "101001100000011110000101101111" , "101001110011011110000011101100" , "101010000110011110000001101000" , "101010011001010101111111100100" , "101010101100000101111101011110" , "101010111110110101111011010111"
, "101011010001010101111001010000" , "101011100011110101110111001000" , "101011110110001101110100111110" , "101100001000011101110010110100" , "101100011010100101110000101001" , "101100101100100101101110011101" , "101100111110100101101100010000" , "101101010000010101101010000010"
);
end a;

